`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
ScnMFhAwM8gXl5aIgnNmJQmh4q8mDPKA3CzwyNCi8ft9rEEbxXIjzbPk96niGlX7U8jytKj4759O
eH/F27Yqag==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UY3JUdvgvpgldhhvjjD7nqO6GyqqeKsaUdn9o6t3I8NaKrNwDt5hxI1QEa4GFUIL3HbEG8tJHdYj
ciNvYB5zFw6lfzAFBpzqRSRMK430IBReUL0+2/oNRe6rnKVHL6goKVdpJqM/YqwLsiYoFXu0bzmT
6liT3CU/pIzx4c4cFPU=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mWLg5uMXJMKh4P3M0iSPR42oFcen2AZ6MvtCg2P4VyXNkhUgggfN6zPc26wdfBQgUfKiu4xpjfTj
okidVaEGkJcEEHZr//aGeEmnh7gFS28M8Zv2Iy4iIZ7gOyyWqL2D7wPplFp/dlg3iHAorYE6+K7n
AeGEqcPYRWUdBrwppD0kodx06rqx03oCAgky/bKLnXW97rodsxpAhpu3BboK5Mq556K1GgfQ6z8X
frRSSbXSP7VaxdJ1C6viU1r+eN5ySj1eElAiNf3jF8ZXEinbSh5cBSoMFKIjwOyXk+fDc2pntzyu
K9gd6f99EfeFu7fPmeCvb7U2baea3S+64oC/2A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eHcNo3fdAJRvnm5zk7oWDFvP2GUQolQ/PIrxTVHyItMfgIE2zpbbMbqEFQkd64jEJiQy4BBPOQTD
gdrfq32OrqajoBdQk12BENQ8DgXlFaKqXP8OWawqKtR2ldKqcmg2vON1J1lmAcvVn3DsGvdlZ6uR
mB2M0S/hSF5K18QwVKDea5Ti3wskfgXH1/U9HEUiyN9ijbIchrxZ9lO6Uo9zq+jH1RnrvAXsbYpk
FGHc3svtQ4ujKu+tNHEdRyO9q2wNfmuU/1rqDMVOfC8/UP8dBo5HjRiNsZSncutMPgp/C3WTsvKF
u9s60b9ZE9p5v2vLmmSSfg+RD6nosB1baUgp4Q==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
JnaNcQiNxMGvvokmewdN4VXhoRiB6Hb6h7KlTM7I4iOdBhMFBbIHUWQSmBb5PmVoPX8xqmclGgHk
FUwKbq+1tU0cp3Ey1hloAULOd6PKQP8qKulSALDa3KSj6ktQnnw4dvf10KYONW+gDCK3Xjaztqzc
kcausTZkIUfuxYlFa9CvPlkZiCRVFch9bpPiKgtfOnkIlxwyRJABhTlgQgUCQdHp417w7J+o+lQr
QP1OvY2LlrPV1j+T+M2ZTmcm4+lifiZlYmWSJWj6KB8VxBUy2LTdP0CZHlYgCLa2M5YuY9ASMNG2
CcxEs86BObBnufKX02nMSPNemq/5xnBi4mkWoA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YZTpTCmEg2/Vx+c9xOJKZs85dFc1nXC7rnhCFg5QbDbWYlCpxOnKebgaRS6EqRI84IbfZ7qz0Wlu
uspcPxX5qfZKPBFoPRwrM3kl9yITeTXO4o4lAkcVtWjB1X1MtRRoo/j5EyYBKzyZm1gb7SxcYQdg
HTS4aWuKnhZuNDH8DA8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jv/JG67O9o7bV/Rax9YxTuprRCB1xE4n9NbrmAmCVvVkI/zmkUHSw6ejOUuGqEeVT18omX8LhgMK
cAFDYCvSdXuuIjbZ7vpjUAJSwuPclC2IL8CKe5quY3A1yTSeqN2ws5C9JrH5nxfwnleoMO3W+RRG
eto2g/6ZYBs1TrJdhXCShplLHTKLXCN9th0XAJqb2ssQ7MlOgGiu2bYGrkoWnBGOHdhHJo9DRq++
0aHFHLLJ6qlxDrBygM3xaRvOFmnMoK/Qjmdw2nCGlIURxwlbupB+/2MxAt4V/EdsybMpQNtWP5lp
5SIi5zb/1+173yCob8kj+GiV5sjbDny4XAuFqw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 151824)
`pragma protect data_block
yh5D+ZjJMT3Dq70RzLE6HHGIvB9QyKeumkX+cqva550jI9y7Iel2lYfFHP2XxTZ4tv+nbfb8403z
pposnvlkTsHCEe5mCObzJayicKSqr9sigErUTFGoS6FhsPujBY/a9QvEwmQdsfeAdt+/Puta5h1J
lH/J9DJH6CJs/C8w7d7UxPo0jeHmgZy9oR12Etybp04sfl+3Vqn1rVDjL7LLlWuBMY3osZN58Kkc
USJ3DdQl989ZQLq0f47qTyA00sY4+Fja0IFrCH1krPwzP5IaWmACZkwFbOdB5AOhDyPOaU93WOZW
D/TiVEUbVb9vqaGeomBdsTpNqPAqm7Oys2gD6TVINQCe/XzuLqwEnylBwY7PYVErJbjdvtcjxy1K
YR0KAsZohu+RxR8g9U5cCh9h+Mp8gLFq4bdhHR5RrqT02Q7hys83LWoMaa6B5nYGlUL9mkuSTHVO
R2BbY1WNmCd21a8LQVXnbYQ+NNGQQr+atDO4/KtsEoEMIjOQJvs2W363ONV/zeda/GdUu3CR2m/D
ZOqznm9AIchqARiim4Jk91qzALDM+pb4d3Ro+RkFLa/98qaSgATIejmjXiEdU6HpoVQsQCx3mUbP
boXEitRj9nB7/vYd0Q07KN5sar0iqqvonN3T47bI07uFRUFRKH+vCBp1dNkg2Ev++jvtZqT4uJ85
3M152umDomaGp+oRK1nopRUvCLZfJ+SzpJCpmBUTnb4f4ZPLhKi0ydmzpDSBULJ76tY1xB7OCtri
W3jpexgEq0lQVL/S5GzydGPn2+9udMiEf2+Cp1+YsvM/CYb5zoaoMEaQmzxVIShkdMApDvEmtCi0
7cL0iyTId6jEGnwS91q6jnaPtaiVmjcYku5Olfa5bnutORMXbfqooaBscI6auW8TK0h2R3g6Nggq
JTyJL4gkYhcd7u+5IrY25kTsNVLenSUaQC2775ZwLbwHqsGM1aKsEc0r4pFTkHAgaRs9c1gbljga
M6UeF58PmfaAiNm7kEoRDhdKNa9AG8ce+CKSGT9i3yqUyy99e5ZtVuZlAUXyFfJ4FD55tSaf/5R8
RaQx/HUNcbTH6INvVl6cERIBP7nDRod+YXIb1JY/0mlzfHZ/CeD5bzl8DnN2CW1z9w+moWa6J9n/
Paqodw8tbyklOND/430vjTkYsdKAA0x9TffSaIO8+rpocg557U6VqhIMChuB7I+bPPhcS8mHUVeO
jqmFe6Vgo9cj4jNF71OWA0zRHHEuhAFetFhEJzOJZAOp5HgRXaXfbvjBtYXAy5WxmdZxChwA/kAD
f+3yUAD6KXH4hYRzdFWP5/n3JtO/XC45z2aiHC/lAN4hq0W/RAT1c13UqRb3zLiz1sYpYUuMStcM
mfOXOBrIv4gC4hhs8s5FxR5dP1VperHPvrAVHV7nNRK+/wCX/bLZfiC/IyzU61w08BWObiahLCuh
MS/7CZAms8vCB5eZwoCMo+pjA/Sr2Feco4F0zibMTg74eww0FxEgzqzYyjoAQJ+uI+M3OyuzPV++
awvwKi5E8nrdZcLm3/JN2mRXf/9fBxYUUq/rRHZ56gcVyJVwn+V2gZboq14UoiyIOBWTf2xSHCHj
YUs88GPYFV4aHnEy9rmKS2W2KngdQ2f2ijzTtlFhVu9lmRkbmPi0ElMMRCIh3Yy7mHWgWENBPUbO
bX4PRTR/8hPk1X9IhXxMgP/1lzG0vGpah/g5yX2oRSh/gZclR0IVmzU8i+3Ej6Dx0Jw50E7pmDIB
roYGpa2J6bA1BBDCeNQcSt+Flawbe1djkhcCbzuvoqex8efMgiDYJfyv59xPRpikbe6iDcYYIqa+
xuorsR0pCihOSeodIXGjZW5fCDiCcKIf27OpVuCAVKrUVaITH+6j6NzvY8Gu0hXp2UTZb2LYAUap
cZGbLq1Ui1ggH1CvNsUc8nW/AGmL2vJ9vfSJdKTQy6wdUDB/DFOnwBE/JUpbUX4rev7kmGaXenLj
3t1i3CUGc+38h6ahDKV4dWdnkVIii4Zhfefh32y9LzdfKjzXDEs2A7a7wtOfTmDhx6WhAaaWdNTU
WHSXx46STH/BFj93G9e0yO374+GXsZHKIJymKuKnr/Nd6WcYj4+MFeTgHjyxQ741QPrjRBnqQrJq
77fELeu1/2LMP/126hvMhhEmXMvMzj00PR3IQifdEx1oWFjXf+ubH2M17pyVfAc+tEwSHizfwHpY
1Af3iHNj+k/EqL0LQuyn0yWj3qXQLzhEblb7K5xJJ5i24mzTj2jyXl8yvf7IoHnlmTBXUZx7YlCd
qBdyqgvkayE+OvSuwDqgc1HrpcZcnl6J5CleluJ/IolVAO6z2sGkrbY764sZ59RznUs9iqUigHYl
zD3FK6p0uMB01xUYt6bQAe7/Yq3VPVmm4Ai5nQo7FSy+lNh4K9Zw9LNvmOC1tJx/zj/hOrLnBkpa
nU0Q952NA3U8C1LyF5KRzzlBb8S6Nj+Dl5GlXNS17t/LUpKW6pI/8jZKL8Pi1mWa9++freQ1faHC
zvCJF6262TFhW/BVJlDdi7/g++VGDenwl5bg4YaXHYOXmMQpVOxdZwoNMv3QukPkoWAP36aYSrIJ
QzyDoCsQJsfHuiJGBrzPCu7ur6EnhiQX/aMRdlg6BaHcGfC+UD8pbu/W5zh79ETZmzA3QLp+i6yo
hmzLge18W4J70t1NLTDuQN6K09vb/nNrUdkEQidREMwWO2xWArv3zhYqZ3oNRKjWKT2J5xUnb7uF
QYoEaAHnfQbRFQJ0mOQn0OJhy5LyMlj105Djfosz18OMoYDZ7iw0J+oOEyLXIU4DKbkLmOzHDtf9
eHrEh6V6jdsVyeD8jO1SapG3Ivo66WzMGsObljGO0lqS2zzDcOdGcB635n5dZEHrbPLku14a1biI
N/UjFqJbNnkOmeCpeu5i9p88ALAtGEpH5b6G8sw/S1DuEEg6/OllfAyOSaCj7VbMRZ5FSnRSsaai
NvU4EYimG8lDhShhSX5VjfJVmWzdY90U3b6a8oZUQTFXH0VDYbao2T9jBEkjksjJ6SP9D80oRq+g
b6HScuNSpO9RUQNcef94W1+tpN7Hwg0c06liDioD9hCQGqEvsJaroxbW9EA7U/1UKPzwYni6mCuZ
tl3rgutw7KcOFNH3ftCLrHYW7QLhwSC8oT4OIoy7YMa78z8eY0BCtIO11vGQ+wzKPtj7p8bVY/K2
3fBjONjupWk4ACwdR9LSodcNtMCjh8UMcqgj4IKa6r5lqIkH3L/FU5ta794gR6beLW2f7amvbQ4I
rhAYPSWlOcuBfIT7qb4QomLsu7sO/FyUszRpcbNUIfXjb0z+7XwWlJdLETQEKezjoMoiRYzPch7m
3t8KRn7Z5DEFPlAFshGwAuDiyq/7+JauWwP6N1VrTpOxrmj6m0xna1oNt86K/Gxsyr2+D9ZnYL4v
zJsaUbet0Q/7IF/GUOkylmOkjAZF8dVXJOk66u9EljvXnFE4sZFXVgnzfg6yMdzrfa7rkDae0Byu
LhjIoIL0y7W6dqZbb7AHvSBnThBKPgQxzvuItg3rZ0Ue1IV1Sj3uz4N7Jjlub4iqN7JyH08tZLba
XJjwwfrWd1LIzA2vR1Iswk+CefPxwQBF/SGXmpErF9VsGF7Lb6ws8doj7Yi3j9Ap8SSWUFasvDVx
/tSKU6SpdOu8OltwWV7FYG996FPt7oMBDEtF6gHlTFY44dhNVYrElJ2IfFjuJ5RDxr9A18/EUnlg
8univR/KdzqYYQKbVyvkCeYcxZ/4EAMrUk3AhABkpsNqh85ulsLr0ln4gI/au6+nNlkpm8f4IMFk
tdDofVdx9bc1ITs4H51Ql3Upglgwq5sgEVtgYxW/mtLPjgDo4whhisH++T5aPbck8maJqfXrJzY3
j2D98OAc1yhNno/EtKJmctWCIJ+mQu9TbMUsBXQ3q0xp2UpHT2QkPpoRVXw4jwneuoDsFuT+jnGT
/a2Zq5Wt/aQY5vHWEnwv59QCg78oFmim4kaJbGdA/KyAI9zbC9zCfi9291pae+QawZO1gJbxMhAr
3R0/bCGlaxklVPdC70/EzFf8Yw8P8os227lBCRMPgKXowlm84BXQDoKCICGMzfG4Tl7Co15TOp0i
2cdC46uOtCIGGw2hVLHXjbGFfPZVflv6l/D4d/wXn4U1diJnnv6Dus038u33vWGy5bXKIdMCl8bW
uwme5DCQYG5kuZsq+psQ1ZgR7Tz1DjUsKCms0L5yuU2nIDSi0REJpQ5IcGizNOt3ENGC06dmUMU5
YMiVCVyQRi7UTTfVLQ33JsBI91OmC1PhvNxsoeQmQA0Etzu2gW25EjzGqM0K+d3SfSJRItOzcDt1
uD7YTSiB/8AETxiZOC6swXoz1QFELH0x64qkAru905FOO696m/puBCHalJYTK+nr9S7fbKoIl6qA
yY4KUdUE7Lpl3UDDzv/efN7upDD1iFQWWT4fdSxqvOUBu8j7+2RYAVIxMGfjYMLnwwWbK94FazdR
EK8v+RfoAGITzA/TY4BbZ/DJyNUotL98ykCsKhals1wEuaY0hUA2Iix6jWeHhmABSFJhPZ7N5iLW
pLoL3+cB1EQ4bDh5RlG5gFk99Mb5S8mzOt5kcFg+cvoPtOOgJoQO2BErnMVg8VOR9a2rqGDIdF3q
59WyZR6tEogPKlWGvLR/5hF507JTR6k+38RyVVI1qKoBf85v8Xn5QQUbEv7+pULIgPyNO5GWXGSU
2T6dUzmBz7p6EWSgYH2V7gAq+e4UprThdmvCGaxLKOURzHu8td3z2NudyVSILVSxQv68q75uxVaw
Bevcbb8pkeekc9g0LpbAZg+SrtzPydYWm5L6L+4aw3F0EQq2+iywR7Hg97Iw00QKa3VICS6beoEm
oJQT/2KXTAnWN4voLjKKmIKW5FZZlxjh1c1cD71X1QVyaURpu7v30nSShskffeV/Q41/WtNLQTvp
d43GxK7P2V/iwtNnhQudCdTIzqshdCGq7UCLrkltdL0BaOg4mYNMhUITkAwbje2nojBpLGrlT7lU
eK47rQJsbusicFpuO0IP0/bkSIg5gNokcy6RuuYsKzGZQcFPHZGjvj90fJYSCmqtc7rmnOaPPpMg
THL6HZWgF7vjtscWuIqb8RCtjn3GrHVhI9mO6Gedw6Y3XfPZZFBtVdkxsk5LOMrdTVVKFZXHIesB
Ek2kAdEBP4hRu5utxhOlWAKCTTTN5OivmDp54xfqOYySgA63f2AWaoAzXe6S0zglYJu1dmgQ4uAJ
VZHOZuqd72GU+pG1/ORUWJ6FSj6uFXNWfjHOAYJYqfykSph/ePQvmFRKbgeFtTd6/Z5Ouzpsk5YZ
zIofTbhygOpZ17koIFf7+sPxjrE8IB30i9OMkY+jOCA/uh6/mRud0HWYTtPUicN5c5Rl3tcpdw82
IuR0RPR6LkfRByNCh1xwXGgbwqVzMtq7aTbtsoQwsxPKLuj0Mqu1veNe3H8i96CLS+xXrPT8leYu
3ptrjD8DCQpjpveb/FbRliS01cEBuVkw9l9yD3RjW1Eg8DLSeFT+DNZXz2rEika1D5sK2qyAUPaq
b3o07IZ+vIs4WQlbXIyozU3WgP3nJgsfCsqlV8o3G4GN805S70nWNTe3VPLm/aak9AI6YY8b/b2b
lzmphKEf9JDI4bAeoPO0Yl2JATRjLgK9WHrL6dH3CRpQEkpXc16+g+b8fbB2Rrq3QbVgiQwkJSnr
0i80qHZ6NRo1rpp865z8Q3Ds5+sJN5Rj2yybOXSVMtPTd2ArCLsjcDRfvMEYb4PNVKQcFp8h4MB5
6tGCha+1eK7TWXowZd+gEg5sHwNMQykPxr6/RnjnZTHhu+xNyoIFk1m7DL232UBm45sMUBCMWORh
3ZI0K12QjUCPseQABfdJotzvj0f1drYUKSeW5XmV9w0KY0x9iY9IKeVBj3euzZrTmkrALhZpHk1r
Tj9Pva6GLKDMOFU5DzqDFyTzGXI3STXdiPIUMxoeLZ4s8PtWBhA5oZlIBb9GBo9iWLIm6+EgbmCm
FNY7TDOx5VMvwIK+CHf9M3m771Y6U5isR/Inx+cQqR71SRprsAJrcd7cJjXuwo+26Bu5VI0mItrS
6WexGbKQS0hbgspK75bTyQxF1CyfFj/nL8/atZdfaerF6QG2/nxDRGjUqx5zANX7hu37c+gNG4VR
pvkbOLrKpXmxMhh0vEXXnttMSuATyiKxPPkaju2pYvIqMStD54EJ/Pfn87kQDhEs+HQRAbwP9clG
uD5q8qdQ1t+oMdyXdbkKwy67Rd1YhKY0+ASBdlKL4JgAC1jmqsmXl5Oycr+AXSGWigLys5OHz53J
agxdeLcWH/2f2j9Z0wMLshN4U30p3k5J3sn+TARZqeibVfd06OZ6XtNB4dFUKKwidAY4OmMdJJlP
ftmV2pJ1/J4jOUxbFtxlOn2T+KMU7cwb4Z+nSsndJFHWuZMyMi4WCr3SS8Hh3CN3FRTYoBWsaIun
aYRoTtWmCk4PQ0Xu94j37enjABl2emE7itTvErhXtYn4HFoUZYDJV4TFGOdhaz4mujG1xjS2+aQz
OP45+d3VqPEkgPZKcCnUFrUOR7kkcaRBH5F3LW8PLpWktKrAET1uWrJieGqPpgP1gGbyheTOJL+2
0bFsctgYWSqknZnyj3wobS8AKPl3am0lp8G0eoVLgQ43RG9yOk05Jz43zjGL7p12M/HMs6fLUJlt
czpLF7GeR28yg2KSQXAk6SVsTK1Ab9aWnXrzdbGYYl0YrTqefy57hBCrSuGAhjrGHphX3+rrWSyI
4I1CTClJhPGwi2+7KCBcT4+HmUWPAHrE9dKibOiJiZu6a/fYuJwZdiYlBV1nXc5kfqvTg849d2T7
tlhSEnCGbnM3dia/q9eWrAeMFM4Ox0edvzdzoYFnYMiOByg2YVzDKnHzMB++M2pkuXpL2HjwsuJQ
PT9q/Cg+lOAoEZnsQJfiiHzphyHjcTKfvIo7eITuSLis7QQr5zH4J3UhWGhLJ19DiePqxf5iM+tJ
3lHwYfoKJ1JsQOu9HUZQCsuYegLt9FMLAoPhuc0VuGMPqgutYmdzg6HLX1j/KgkaMQ9iar40qH9a
zBe9tutLu+XxDS9HM+KWVZ1QBgjU7D077kYqPLqL8zkjWqQNbEH7vwb5fSFeBSr1HRVQGIIfUrJS
syGBgDypngize7ivntyIHWnacmFrY9M/exaiZ7XPT4Kat6MFBHcCuURxWj28QVlgXhvoNFQWU32L
/iPiK291gCr37fN/2fhmZ0npC+C2z/MOpEwr4u2byo1pSPXe3hE7oFGe17VFhoJ2DJ3T8bgO6n/f
vKw8pk/8C8b2pocIDCnVDn2bWd2JZVc06SdVIY7kTU1e68E1ECaMPxTnQpPD50DCMNDDSGNQ7A1L
ZHQadJJHx1WglUlITSNObjYC281IIXM5dTuyjpDwAzqnstrdGOKO2rqsYRdHV2e0ax0raYg3K6ZG
lXYqtooMcXKB2MlXJC6bSF3zMg9ak93r4qZDRM4yz6YrvR0RZ4jVZ1Tn6mAgyEl29l5VKDpj5jB0
rH8Vq7FE0JDu1+bqa19LUZ/pd8GPYU/dNU7OHjWzC3dFNefiutdW2IKb0tBJ38HKdUKTvMy+cj+2
SQUqCtPALOQtKg/T5jOkFbMBpbQCiijxBb43MhWFSWv7SRJ1Xl5omQ9RiGBom16+qX3g1gcsS6pD
4Rk6JgJOko6F2+yy2T6IgMdGjRNVW9NzZ1s3tQbXki3FJsgGi2rsI3V/BHnbCJ9ptLdUvQPjtO4j
a/V8O/89nfgc6oCybcAMET1/WtPKEPRQ17n3tC1JmI6RYRDqxpMCO2zWdsHoXMhRa/er9NjN0N95
O/epZHbMzOwds0i4XLSfwXTUg+wyVjel2TW5ZI88qpsLXo7YaspEweD99449fu89rDoccwyYEEjc
OBf86tk3MjDJrbLF8rZEb+o/WanRPhAz18WPlNfpGbVh22wJzHYXhAXPluZz6ozJYWM5aCaHdhKy
aTCHE1ht4apYi+9Lfpjv01cd9v2/N0rwT5n+WpSwtbUxVXQTvn8Akzzf3DUsqqYqLuoRgezjlhEH
dwRcWPtY+eAZZQ/P03/ahtBQGaZtwnuiPYHRitflvud6SWGJqSVPAoHpXfG3wA1NMoS5oooqc18e
aYKWyOd+JJlC0KCKc//j318rh6GqtAgbTuHZwX6/loAG5v7qDibsG73YBjOIWM5hudWewi1fVk+R
gSnqJk/o64zTEwnKIXzz/ZMl9pXhLMxs0XbohDLRTFTiidWkkJGpl11PL3yaCeXPf8V23RPFG/d0
khhOTMMwCLMHAibIp/NsEpHMVMzKg0G9fQcRI66BMsMY/CbCnOwoH2K4pjVh8vmW2biXK4nVly0d
YtnLskwooGAKTvCwZyNNGHHI6ZW/My092SN17GZoYlZ5gBBV/Zm/I4yjGYQwiiwMKNn9QJuyFgz7
URklGSNUdf/OpaPywJI1TFO7nHzwLeHtFPemjLrHgfg9R3IZtKiKVopjjLR89N5+YrJOvk4zVHwL
RIEyOphpsRu5J+KeMc0Wqcayeei8GPDYjWGpReTIowwnlvvFcEt8LOD1EUYoqLzBkqoe+hHoccdi
G3+1Z3OprrDy+e6Zmc4l6oRuFJb5A6DfGbspEu+Af/E1jUHzbQEnZ9odVOikqvnFmReV8GXdYZLO
OUp4CnyjB15ptTaAZXiQeo12jw0ja6BU4FR4tIc9FmLDaGJ4uE5OKv8egUaGvRMKFWYBhYH6rO8S
ciXQZRkhrE6HkFpa+BUZjjJ5YhIlY40nRQhmI59ZclEsu0NN5WZsOnpMeQG/G/hwXp8eY5W27SGJ
gWytWvE/mADhxiONGWZKfqoiFZLWeToG1rtSUx98w9yLynwGsFN5YM19wUwmHL2ehU6g5qLFT0yO
8vRzhBSn847wAEvtbtBKYZCqi18Hgkh1VSD99kHUrkVYd07t8YtvMjKw+2nKCl+G/Vz37JRk50xX
OvDS2Zez4NjBrkjyxxRsTzbB7EPkgzdrRou54lomX36ZFnGHZBL3uPzsRR2TnlTx3v4UBfrpBqO4
AseqIqzyV9wFgI1dSW+CliU54cVxwGHGqPFa80Kb0tavRZCdXNQRpDY4uPmdPGGuzrn+PL50lz5W
qd3GoH1Xr4D1cRTCxglxm6fuR4AqP2Xv+fvBlpLsbE5EaQX/t2uZnIUiikFqyBfXWT+MWzfBye7U
CzpAzzy/hHvQHZCg/Burbng/bFUC3005yYI0nlPAmSGWZ6n97KlA50g2zhZpwfv7qdilEJD7AV4l
E00+ATHVVd0oL+7cc+70IBwYmXSGXV1n89mtaZEw7ePzX66lfmZ09Ipq19S/AB+VxADgun9eyEDk
YswSDNfMpO9kz3C3kykVeuJZML18K+YkPd86Rs5jhU3UW/ifc447UyVVrHTgAFvavYCgZhReuAMG
gHby54VARHRUu7CnqGPgBI24xkUdAniZHrWg5HUYSP2K8WU0KtFHkyKGyfZGj8M53uqDMjJXJdzw
mCwefaUSTCRB/yPyQrBfglFN2h5U2VolDYFN3y/wQlIVhiOeS5c6zTQnqT5Fe+6BaRZCrQHPkqy1
q4YxVgGdEIKcywtlk46isMWhDLSRYxmoxleUz4JMhfnMQXkqmda3WW1W2ow0jLGM5RzrqEsDNayo
r4EdzKgwCw1Ww8gYUlBY4/jql8c6nBzmJeVpQ9YC7J2oc33MkpuukRnSioa09q/cyQhxICmr6mKD
FGLPpsKdm114tXyfhIa5rGWAEhmBwQqtRbybR5BtekwCAXhBTNFInSCcluc4kEa9jeGh4KkxOMNE
B5amdxJPo0cUuETn0gU0WldQf8c7G3EzZpAg8rSYas9pcWNf7UQibcnRDs/qmXz9F80AjEW8sLrf
KfqpfddpFOrlq9YKI9byINvgB557fAk51SpwgF1JRLDMKAKNw5B4zB7giVzAHtmnk+V8jq/GHDA7
75KAel4OkVfeWTFDy4EkoJNsOjhhEFHTavepUN77e4XQdUnxoQmUN3T9ysOQ2ca9t8Vu63qkaJ8P
+7IVHh9O+3VuGCdoqqNvrP1U7VsX+EVkXpoEfdw6F6vC0ipGT+NeSPm087hwZvLpKt+T3jn1uszj
lQxW1fnMLaxToCoQbgA2WJ29Pt8zSy3Ahdk6olOrYVl5yOlJqINTuaS0B06A8a81i4V5KMV39xud
dlFNA7J1Yj7yUsOsbOH0D1UEn4xRsCIStKMAPRGjgyf10oQgYyu+TYTVxrUPjD74z03IeBP6T6sJ
ST36kUR3vgIx989IE2F2f/eVqM4EhZUJaCJ4zD3FIxBPJ3mzEl8EOyWvIpDHKGU/GmIR+G28pXbq
0ayEwQzzzY8G4qCMDQ/uA7v2pm8oh1rfcsIaZxHj+rm7kTBaXCMHQuzGerUQ2kNfd/iPGgGAVqzs
wQNxMC0VypgfApcmXxIydM6noSBz6iuXiYpgq1zx+s6FTdr1aArC675igYilKskCWBghplxg0WfC
n5tYKXdbF7FFSCbInY5ltNjUKYdAeUVE02HPakHHFhXBkgvp3gGAdGNfJppl1PlUEjM9zG8izy4p
vQcfX/PonPb/+s3kx0nINSvE42Mns5hBxL79HkSVvbE9bbbwcx3TIKgq20t8EhtFvorYAuEnoUkZ
CQaTciSAs3QRpudlYSMG6sIqfPoQ5nJEjoSgHSEaq9tnoqaMJrntqdLZXx+d5fCMETSHj+dJf1qd
zWE0AAdR4b1LQpnWDZTwTgorCC6xUMU9wWz5rVc7epRj4wgnZPbKOadREL1OLP4TFVcZrgpiruSB
ihPXwu5VxEc8c91HvvivozZgjHdxRxrkVdp03/91I0nGWtSD/0PLInu6M8gCXT3saXcNFd5vvFyv
Q9ABW433tyJctuQT0fCmkrPYT7hSm9mNWStrDz18aAtx4eO3Istli5mrND0IJJR6+fZxBznFlO0d
DeYV1oGalArRdCSMV5ylHOLzoBZn5QtABl64fma9aANYwhQIByy8kZQlu6jbQftwXy9rZKQTXuiL
5DbwkDvPjNlWiABqen+ekO8NZse4MXYdsFoUSp2Gu/ozisFI9lOnaKIgWNDrSkF51/8pQqqIdWEr
IGOIRlMbTqLW/mkTpOJkD5wEiTvmeturNJsGX0wQZ5czhOMK+kTRKuPjpeHROHihJAccm2V69Pvu
BfOjPiQZOSPwHCYE0kwxEtho+IsLOM3Vtp1UbJuwDYjiWLTneQYd2Kz4+tEX9M308GUjPQA34dBP
9NrCVCxrtLlIir1TMH7gqsszapzO1CQusZbAzpHzDkxsqngpC0yVEOsBPPEgs1l2IWC8iSNYg+aw
F5FIZBSt5/bYJSXXZcLKEnKsUE4MINbmCIxg35CV5Sy4cb7URDQ4znl5ha77+xyvFiWKYqymoX0m
hqfML8zMPLv4WeWq+mBiRs6/Y1uF0rM5SmrFafrlfIf73YXMjLuHVrL0CHAUr5t7DT4RPuSPIQVf
4NB9GYOz7OG9TUc83iHOKcxsaN4P4jl7QZcrc+dYD3jo6+KWSy7kt4+PxtdT7Vr7iW1O8QXJ1h1b
BztBRNPmGbDtD98ZxBANkxN4SpQoldQI8q+XfRhaEuqPN74lfy9QBk4u74CcDmv4V1ORpc+MQ6AM
E1rrU4vFPV1xyYFWTGyJQa5fOprin5Sg4rrjDP1wdjm9WUiSkDHPlwyfNIHAUpdhZxF01bh+K5Y9
1r2F/AsCmlfAaw5162BSM5qnVr70v7wvoeAm7FIjgFknlYdcDPFeNk+fdrMlHGKiU/WOnjSBkNDl
9G1e3deBBkkQPKVPMESczGoyR+r5J0KLIRAEHF4WXSVpwaSYu+/HGzs1HlpbURtbfaFGoXGpinpW
Jpp2nhuySesGiR93BeE2OOaIFDaho86SOf7KjmmGN+Q1jzpTvNMCeDxxT7pmcg69UZkWyjsCx+43
7RVgUg0Teji4MJ92a/3TYLDdOcr1M9mODzj+NBIzIRxFOkJNjoLUnzfFRabjftNw/UGeGcmlbR66
H88RqrzPoDgMLVwPW7zFxUiSJRgKMZ6jRKQf+39fj9/piTA64Cq54YNCxKbmifRZKJ++TkrCq1uN
BLqdyqZO+3OXy8wHnGotnJG4gIyUAbK5ZZQID38BFWC9gDwC56P5xyAOgvIVnaJ8uiX4RD8NgNxj
2P4j9qgEAHB5T/QzIc6M1N8Ivj2PMh3lnvIhSiaUAnvvrop+QiQEmfACRvFjCrib6H06TGAAx4eo
j9z8MOY6DpPTc2m+buczTWzUvx7P/uvJp0co6VD/x3ZdImEMG30Qp/5RP/U6kSJ08buF2lfqNhDu
HqzxZIQHgCHUbxWEFbU0HHivSJ8Ph4Mt060pOZLeEO721ZRpjvHJP+MXb5i+//xhlQ9HItZYysdq
oWHat6AEbfPs0iaxEhQC30TdTNV3jd/XGtzgbmDPPujrKO940Fk0DUYbXD8XyC+AqThNoEVxybWE
Vw915wPJgI++WYIeTz2O2sAJYzCWN4W5X16Lbkf3QcMkL4jXIviX/4/BwxnDIt0LO8dsvvX459s9
9KRqXWszh7WvHwq5qCL8jLh4qKWaAPYqOrgbdKO7E2tjLvCKsVqqBGCieXvkcGH2nerGz+qio79r
90o3KeRFVuB8PwJKCdRO+nDZemQ7yb6FR41/u64kNJK3nncVFtCewVJj6Jkqfs7I/jWbusFsArLH
41OjGTU7hb7599bJ3Iyesb0o2xICATnxmyNVsgjwA8/o88uxPJtvbUy0mlxRz+xokL+wCk4RqVHy
nfyvLPIhTVveKRX0uXv4BsUkvb+3K2Br2q+yZao2LmMBptuL7WS1JTDsd/BFwunBMbuGoxAqnvpk
oXIVTuH7ymOL7MxWgj1VTRLv1gbgE6LQ3QV1v2yc29CJaJYP3jOdVoWFrF85Y1cqNJIspI5O7s1M
qW/5ogZTV7e37GKKZflSb9TNgBGdOdzlubTfaHPq+6barNfnwiLRgeTnlrcPrAsSSNZAXjhrw/nx
xVkjgczFiguGUbLcT+HBcUgk0ud1R6ZyL9Rx73xjLWXle30v5SgrC+k42aFkPTZslpysQ0NGNtVh
lO9faaFWHxfy2c3slzfseZVEagrooyEwRqycYUh+ZaijB/D8OXGl4xMnrktOtLY9zq9I/qMuDRvf
dWx1gMRtWcB7/djexVLt7CiE2RiIysax2zhp+mRBpRCCgbND1003gG2oiaVJXvHo4XRgANqXbo3v
kbfjOd0SnvkVFmexy/c8o9pMfjAQtw37qUkJ90sIvP88iUqsWNgieJdnRl6gb/tu1d8/fEJ9A4zG
mMIGSeRiYOD944SC/9CP/QE75+M5JA4fctOO93ZlVmBz8N1iZmt1BohXZFCQbkAnQyMw41flYSL0
OufXFENIfIznn0cYWV2a87xECWtHnFpSPYmqgv+rPXH1NgSMsvKLgRYDoCH9EejP5Un0EjORWpKN
s2U92Mt0LDocDgN+uuoU+vD5Wem3m0yAuHWQ7yWzlGYrmacvUDjafRUiEPRV7q4f5AmhdIO3mCGR
+hazzE3VCsLCqvX/Wc9zIzd27fnfcvw/VwvJ1MG3ADQL1WK9gJi4i8YBskHO7N95UVHXKSVA9GAp
4/T4DIoojvSCp+9pZgOrX7twcV912+Qg7D8iJdlXV3MQcHwPTXy1KgZKO8Tk8hb2eid88zyQKirv
ANFAiMOOtkik1fbEqs9K1TnYSy6SoSCB8Svy6c0kMKaWcCOaxHYeD6oBzEUhvM4VBk3Zr4x3F2bk
VeYK/4mTDsOnsoiutX1W+42BxrzAw5oUi2zR8KLPn3fgDIKa9iMD3iRpzOSPkK6f2PHhY5vSZhSo
NbA8Aaz2zDtyOHsScoy0DchbFfw1bFROWvo2l5MEVmXL+aTwbOisFjx3qwCeLDdeC1kYLo3OU5bP
1dccmDNYimeiID9CyYTqwpWMMiqWvy0K870Lb7IJFya1uNW4h8DR7eCgYAdGu6ESBA6sdOnFhlAW
31GXw4kYYHiFYZ3DA7XG9PGW6kgO1Qwij8atPrnp+iNpSuVxgzY8LSyYrG7x+QO3JvKjwVey5q5k
xz/dYdKDl4IYj05ub9apzNm2UJxNUTe8nlv7diDJvHGEtwT+msjzkcQcCFM29swGL4xDS94lAY9Q
EJToO1P9VoWLghVhKnCLmeoKRRuoUuDkrDEn4D2J6o0t8o0mzE897PWUJLv8K0bMLRk58VC0YGXp
wneFPkh6VJxMbXRkIlgt0bauurzaLtv74jIMRjBwFtfKlEA8gk7+TJxFSsN/uVn+Sh1i+6blDlFQ
IwCHzLDUpXaK5cWs8csTtiSrZPRuf3l7hZaTIcdbMvkd58Dl5tPx0pPQQ99x5VEBngk6SkDYuF7Q
EaO7jWeI6D8d9dmP41LMbijmT5PEuzsczeMwPGfeOt71b4k8zsDVoy0EveCAGKDQoC8dpTQDCplz
og8MIfz1JaxKmryi21n7VtuQJ+KYtHpBLrsXzSUwWVEMmVqFixXJjES0dKx/g8tTVH7ofA6Pgaoz
nwXhl/TNTM/aPWkBgyOOWEnoeDURZ3jCJimBzogOhpiwG4hBb5Ubhukgmvsp6xYgC1PmzQmM/93J
3nMx3ISq/5A0I07yfRRbcLM5DOiUUD5LrZ2h49KcIYSJaYd+9DMp/2UAQi9uyFv1877FfqaM6mda
pESmKGRuS4pzAz686miGvCWA51WuReeaX/NuHwP/WDScXD4NQPFQ7WkPjK7VVRKGwgK2n7pZyL86
wqjUQNwohLrSihK6atolY4tyklRGGRhNNZhOJA+skkNWl9pK5f6x3l0DCc9gzCrzXi4A8OfhRWUz
YkSfNk5sP/SAhCJG0AvoeWzN3ZQ4DEpPzEqyyhr75nPfhKehvT+Vd2YDE7Y/xB6jHFIOLIy8K0W1
sPHBVp8jDQMYiwTWeEZ92mWrYUMtY8Mx5DPyhq1ImNYZxKCcPZ23v6wxjX1eqMr8dTQoQwb4ab94
JI9a++xBGlXGBPWTql5qYPaEgnWPa6tovTI+qjxIt77aapMW0qQL+Agxg4xOWCWImcGnCVYKniMG
RUDkGrwoayuBjU2GbG0cDTezfs5W9Q9w0PXDjtTEpT1Y7odGYGJBfy15kx3TDi7WMYPUT1T+25Fz
rlcb4hI0E/yxXOhrq0V2C0vhS5Hzl3KjvJp2lF8dt0O8cLzsejdYT/QOXsobp8AL3CibN+4PxDEe
6q6FVXn4vYi5L5iHKx928nqi0iNW22zAeLQJhFzinkfHm4jSwJUO5vESl540q/W6tu6FSowvRprs
WWeuQcBz/27a3f2oUJR+yBEMKtEUcCmxC8YsKBemvdr8hVerV1+nQdt/CCnPWqLz93MUMkh2vlGz
xu//f6aW30Egb5oWJQ2/IEryJYzjBp/FezvwTY/3u+06si2zUaLl7WdfvnlsU0mPIecunTZ5sVRG
LgoTuc67MH7ERTt5tNsjtMvCyi1AzAtwy00H7PsNdtlthjJhouI8jSkCfVMRGO8BrPU3zG4P6I09
07/4tujhVzMwit/oTa4mHeN3uAeYf1hEWdhZdPcYtESQuXX7lG/zjlccuGoJSvR8npUmioIJTfjZ
9mXkvAoCULmjoHAQju5h7A0N2fYp7h4rWXxcESPZsaGlt2v1EwBTo2gCInWFka1ZHydWKeYzO9jX
G6uUlOMWr13sKGcxkkHcHT11z2OsxRWERR2rpUo+AdSfFQrGfylZ0cPityZ5wjuMfypaz7IRO3qd
XnAdEKe1xsnA5t+kLPzHNuCZWGlVLwLxmxZ4lWit7L4DaGZIbEKuPbyAgqtvK5oIHZrfgM7PYP+p
7R+4R91rM4zhkZTnzT/fNBLNZo1TgJ+9ZS2E4xbCqXFg5xb6JSvJOafkbs3W0YonSV+/g5JAOwa/
Rz8aPmk64XBPj5yqRYf9Zdc7LV4+cEbyw6MN5dmDGeGbbDm0yolqYxmCrzHa3ZTQFsJ7EHFM3dyh
PjYeFncBRWiAh+90TsQc8YeBRObVuKanzt6ha5IiburYiDEnL7XtXBH5eQDO40SlOcjcZp5labZy
nTPOe7DFUuy8jY4UBpJB2Dlf7xkNBtV0UmVtaS5q33wcfqHOeZt2BCJdS8+D0n+a9Jp1I7stYBDF
O4w6wBV7OqTO6eUHXlMZRDoHC7yyGw9Q5hMbWC5MgxEyvMbaRay+j7aL4hZUyFXMIKsqj4a2enuA
rE/gyu1nFyai1orAVuBZgroBhaG1b6TEsIJwzAeAbYjKRHdFpG6Vv5X+ecxnU3aKYezg5UHDc8/u
1M5+CZ918Ye93LoiQxEjyNVZEbEVItItkfcyglWKJqHI8bQfIVCQ4yraG1xxqCX2cUPPLj2y15VB
pZtm9PDrHdR4NHZFN/aQhpdeLZxpAz2Wxu6ZRU72dV5n7KytrlGQ3froj4wFuVSExgfhVHcRnZaD
IQKZKZmjJ6nzaiHw7A5v4LTCk9WTkTiusT3jfvbmCpInXX3wAgKUPshZ+yaEKI0/3xspDH/Gkw8n
6VDqQ6AHm8BwHwy84L18AEiwKTqhxkjDDQ+pzQMfAkvCTSsvDV9w53h/+CrAUDJIw7b5nXBlaNEA
UMfSAIIaWfG6BK3Yb92o/51wYdu+tR1ws9dvwDMmr/SrLcQpT4CLECUuQPkPHcLaeBl8BKSfEav/
HBlxMg3pB2Qt6uDjbiXFPLiIJyoeJoOynV/mNslOT9PTEW3Py74HaWp8RAuZCOR6SmhXLTR4pE10
lDRkdsB9RbxhPRV16MnxYaijFHBSdjJtuLp9kJlxMmSex5d6f5/DrTl9kX9hKZGTGMI+xUJxOZFS
6JkPGsZTDv7wIfKZ14MlieySC91h+RIrw5NSrrlRkM4/grRgKMqjJ34775IJjNyfN0l0uenaESu7
ndGGtq8MyF/76ucZHqGI5eh7qG7OMomI1iZitbNv0OgTetfVFztTWW8QDgf7ZO4Xav/CgCwnUR9q
k1E0COub46QXP4omkuY73SqOccQdrKX2jz/SDdSvpcxEtXO0iaPT8RHSygEh0CExA794A5S9QpHs
Qg9Z7XhSct+Cd/780GLjy2lLnyfsSVSjSl3FvJ91dlwCeMUhTeGeJ17gEsA8+ai4qU9huzOcH5N/
1TQZq3hbfMiEkDSGJSy5oLdWjPqHrjKLOByg1bXxlZ/qCHnRYzPVYiFOBIfSpXglKGYCS+ZgdybU
zRyknDZ+TkysM6CkJ3Kkj6UGtVAjQjOVcwm9utxz5Qc/+0wMhL6wCdccQ9/gUQmKl/yTgoPnzCYQ
w6n0Q4n1p/xZqMoJRuG2hKLkzwKASOLtYCmiOKW0wLrVofgWYQvePJxIrFNkiYVdvnBJgO9eJNO4
qaIC24ogBDDukCeUhLJquQc88MiuQDkP0W4BmY9eFlxv7NI6eYTXouKSD/WdVyLTTxKSfZvKJkCP
4QuJLwW3JgO+BnUGf41vZV0Viloq4dcf8mSa89u+oOtZ/Pj765ur2xXONDVXaCWkTxSslbs2YCAZ
eJ/nLeIwZn2i3CT7GBY/MXT/it6dXyqhctMHplWsImb0Vkr8+wckelf8olw1Mmhsxkerw5Y20FG+
mvbMeMvhETNv/gTrbk3+YjFOnHipCiCA7iImuPm36NH2u2IKgrWUevAMue6SidBOki3v6zWasrRl
eKL85t6DZ7XDK/Z/33CurjhDd+hwfXiQ5bp5z3KQZyJoczD0x6Wa1uS5v46XWsbhRlNqZQvjzSbC
47wNcYGBWUm7PqYTEr9s0iPBBltGGBV0is7fcG75cANv8HrVM7ryvsJG+fJzGarkfFsFpTaPlnA2
M2gfVmpfDXNyOHQKIge8mxp0gWTzxhlkzWpRuB49C1Llj45hKh8vQB5yS7a8mvej44a8nS0oR91G
9Du1zOUDjwTIO4NsliThRXgDoeqyiFtyZBmI6ay6gZ2oRU+weZcT4uTEe81uyX8NNQZ78A24HtGw
R5WdUw9LVSMSdYYMnS5KxOs0NrWLB/0FTp6bWTD4ydkFCU0xC8i+jl5wDYARzCtbW6/Np4EjwVVG
G6JIdKlpMrG21T0flz9bY2oBvizYSqkXIDoTMykFkX3Ps7NwSItq62nC0/8qVcFgtuGjC1Vmccwn
Mss7QNzPe5WzxOJoT5T+Fb9SkyGevE6p5ZoNypeKF8Qd1iiieBf6eLmCLeV5+nAaYeCT+/OmB8MR
b1cBntwCz6OeJXw9hfbI2Dq7hwZpG5vz+AOyt7bpToF8uVNhgpqmG6/n7v5xNjDwOiJd2i0Pz8VE
vs9GL4gAKsho0eatFTAdjOiKYiRk/ipy3Hm4UOLWCPAuMPmmevURy9vuMVJA/UJoA4egS5AVS+pX
LYOVzy8ZBftkmwO+CDTtK0XAITtNsOb+vmEWeEtbWQjW3hpE6C2kM6PZJ8oqqx9YWtDTZ/0sg2NF
9Yh5UOk74LdcXY3uIVttGCEO2KFE0moqDlJ7nJ9QK1l71TBIeG1U72P5mYXDT/OPJZDhsh5dMa6f
fP5XkLx5DEAAKG13RnWNofF/dZ3R1cErsjcYfXrcWtBxibBtbZVnd15h8pWCHJWGxBygniLqZ3nS
B0LOS22jRb+0i8fOSOSP9rZYWHPOESdlXLXoxSCVoMvR/9yRsfjq+rvq4+wnsIkbpz1MolV66sMa
YQqx5FKUKIY2hTRBKuMIPd3Gko5pzEw5lQc3NiUv45t1DiGb3Y8vhXwJaVAGf02SDS0b4KRO5OX7
sVV4s4meFycEW/qmlmViYHHdOoLQBdJmo/Q0Xy5XbXGTuUMcZ6DWxzVZCIHR2he8YAYwL5VJLpRq
fFAEz/qJYouVby3VmRTukkutdXWEK8e5W9Mg8EhrmLAIFkdba+xHGD4q1WcveZPqLrV7HI0ALGDX
6m89Wo6MnBHXSLF+9HIkob02iIp8yVQzWJ5xsCGf0Pcm7o4nsRsdC6pkMIHHHZWaXzqgIbQOxF5u
qJBk+AXCa43hbGtWVLsE6LJCQPpfgAsUvKGBmypbG5zyLYYzaUYUBlAresE6aNjjPp0XMjD7A+xn
Sl3bpeNREuGk0gt72DbJQZrePSdm/LL1G2S8f44rP9ETJUU8sZSygHmyXUuWEu2eYK9+jnY8PSSi
joz8cCLrYfGI8/xxPQMyPCCh9aDq+ul7p4qB64E9aEsAgl5Nt4kkXD0kTKbU0VspXPLe8FH3Aq8R
kXx9tUaYGyhWfzSzuFfoCudhZD9vTnDITRIJBXbDnaxPbocW7FHWVYWtnvTWEChKhb7h3rIz7LnS
oNVrwiSdlCfhjEyoVnuEUZBk+oPLbYrJ52jaYwb4apgNBMElGHdwyOaLxsANDiaFtZnnEon2BLei
h500wgNbPeWe7DZsa8ERVqJWz7fe5tLl4Z8+ODgfZOQz1LRP5UlracBCQsx41X0BCjIjLWN3Jf5M
BSNczPvoj4/oKXW8y+FlE6rDz4jtKSxMB1kq7rPZKMpt2FFJtclKGZ8PLrUN9aSFHJ8RAm/8Pu2R
ITW4SBC5D9qI93VWkKahx69E/Lv2biezYy586G6fWtDZvGxEu/UOPzeS2Cw4iJOSufHTuTBMJKh/
WsaSwqQzaJwqrQb4KuZVjkcyfhtzK0JZf4lOrQUSzWGLa8GZMS1hrxRwvk/pngjiOph+mied0c7P
oXPo6X4zI6W8Ax6Ts4Bs1kK/d+nCeTAHY6Y76kQ/8+48gYYz0Zy6QQEN2V1+ppYNNpSroTdibJHD
pk0uWw7ew0nRaeXLPoGYtYNItT41Jf/flC9LjNVa+lDMOJmGD1acxhBvfyVa+NiOJInhq4w1rGdR
5JNPiawKGoufcLsjoRhRZIwofhAKdfIgbx29ZMjF8rVAL8vSjF9vm/2pkKgkK8Ah3ZPpi6PVoqgB
5KYlZT2PxdiuFvSXFsNODXbtcqSAnP/2ngQzSl2xKQxL/nk5XXzWYEm4X52CVP5qqQuvG9qmh+hb
Z5HyY3o6pveTHnolXt/cSWdLEug/an5T2IVoG9GnEuqVQ3BYBz2jSboq8+49nhTohBd8Pt5TlWcE
fzZ/R3WK4Vf22HczUumf3Q4VfE9950M08s8hCzV0omEXxIfwigV2cNCfrTMAJOaEhCYysHjAw4FT
Qvl9J+EHKupAoPQ70svQJ+4V0B82Py8Rk8eMWzeXKTRos1GVEdWW7H7C7XKH1a82dfGsvwnEHi4C
Mzk8uvo8bNBlWTYy8ENRkUicIIFbiAVWzNq+g1bMn8Ij4Akul6PeqbG7OeYrpH9dyBr6AgCMDy6A
/OcXNW/f1Omq3bv/MVLOMRMvQ3OeVlbQsTTDLXMpl4jbPaHJgsl6akkSkJN2KSqv7BQK+xbdbxwe
XI2X+r9jZATCRdQxPKH+fghu1XN4a7g5MYby7uq7o8pEMliwHZHwE1pEFtAZVHY6Evo+i2VSZvtW
pMSVNj0D7KKFfCU4UCzAjtWbgH6du9Em5uoCJhjZbbMZMC+YZCzyFJ8kZF5/aZF9BA/c4dZPBWvh
XkNblbMVWu1wxrdVSHCQ9MMOzyuybqrHW+LRLoSh/eorpRwKgWEZXrLV/OEdESMytMPBbOL+Tnpi
ihHWk3Q50uzqkJKuBOx+k7KaRpRML8MUymH7J60tzHSoIe81vr8WNvs+Gc3GNNnUZFjig5+tZhLi
0QDTuvIgGw7sYfBGwyikAXfIK6gZ6YOuDfh//lxu2Q0lWa9q7WE35W6YLCHU0GooOBwDsWenzlM3
pBallxabM378OQINEGxbzOZmL50kYKEPD0t5Hq6SVTO2l/WI6NsgMSET7tMgS2eukpzzpBiCXwuu
LnJzVUreK85FeSqvkDCt+tRlt0AX9rSyFZvWaGTFUH2FMvemKXpkV7DEBsJ5JnI4BBcl4JifBcZK
1SUxzGPFgu4cUzGVjwfg0x7J7TSlkgSEVQJzbi602xywox2gs0ibwToKgcGbNdDSws+nM32QzfiQ
7lkvEr03M0vQsXhNzB3S+UIhl7fJYege2jPReRwauPc+EYwnuIs9lc3ecRsGX+MptYdH4ZyWeKkE
YPs27fhU9+ODsY5h9W/FQcxc2FdKPeC+DRAWlVR79FmQScoRYbFz74UDFQ5a9BKwt0Ea/0Jlr21c
bd6CYY4qeoSCo/GO+Xq5qUvZUkgwEpn0R/XMCQlj9v7YQXdrbWml3opQ1qlhgFrnPoQHiddUjG01
BGTmsOGILHct639yEhOvapdKsfcJO6doNMs+JnCww1rTGJvF1iq/mT4ftrIuMqv6BRQ3AyIIbE9n
oKz47NoY3cmJehUbe+erEkhBUcQ8R1Q2pPjEcjbA9HHYGtc4N8bWQpNrKNfhKXLLNPkvyHvvpHUp
Lzgc0/krzB3FPNa5Z9bCYN5er30TgaUZ/tTAiQP5D6Lz4GC0MNfY+m1iCs4g/nTB58YlQUrmpSHs
q+lOToe4Xl6abuwPWtaEVoWMvrVLqPVaK9edVfhNlcSdp89TBuQjt0kzg/sGQaMQ0TSdaRe3+iDe
kNa3s7f/6WKlIsYLGDZ3Q1ELvlL0zM6TFZM0BxSR3+INyjhhu8tt/k7hUCQ1LTtmwhsvCXTocrIf
qqfdhGbY5oBvWkYnGL6Su/4vt2ORXTiTuEn/I0/JkoFiIZpHVKfkKUvgeLk/BsjPytVDQSA19yur
RjWOHvkMcG8J0egOwhbiZLsLCuNdAG8VIrDxYKC3EsDsL2fNS/Gcldogbg3pQlB0AmTgCeJrZ9Sr
2duUarIhZ38axK8nKI/Sh7fgBIu4F2u8z/xrjrIbuIm+M6G0X910M49hDJzvbBYWKTy1K69MCmIj
qYGHv/mkZyMVWzFzf9cQLMhfLllE9ZSv0YFF1Km77M1nXply2H3nchrgB5wEtB5nieizfIa15rbp
9K8xYe35/d5bMXuev+XyfgNX51thIyKlE2zlbnE7n/i0oP3foP3tOZqVE1C+sZXW58MkOq9VPUmA
rhI6dPvOw+XxGS9kcyjdFNXtkPrUzyo1PIFqgHtfEeG+WoJqz11Arcmqhvpx6OyuA+KHnh8H2+sv
gU31mVkuapJfwmntoIheMhrZY3Mcto/X0ONvUkLgI+nWBm2NJqUOkph4+VWOOeAqHDaPROs+0TQg
YvAUz1M7oiapVvwder1ZhFxZItGCIn4WZjgL6TAMhP4ax6s0Fl1gqlEd7+3V1QAOzwzblHsqqSuC
f1kTRs548ZqTNZ1aLBFzRnr/eK7Y3NCcVyHU1QiYuk+ysDFQ15kKxUZTh033eg5k8VBysGd0etKw
YsVnJGgoaTyDa9xfA2cr3CVAE3TVYZeYnbKptCANxiTnKo7dRyB2exQ1fFIOIQVtsX1cDeELAquK
ZLzWu5N/bUXszU55sD+5VPZS6H9Ik9wMCvymquXMYTeYUIiEwMFQdMncB4yc1aHcJQQFZBKl4lIV
W8Prx2ETQZDzpCmzTlJe0SIwYarPMfmMhIWgG4NmVn22X2sbvURGaLbanm5OHkle5CtPHYtwiAgC
TUYfCHyN3UxPGbNkJ5V0taEFBfsw/pSgpthmgOIyS/hzXDceA3D78TLHoU7FzJXjfMD0K5+T5FKG
BRvAYnvN8cD0AlrEYqULb0eJGCN2Mge5ARUw5yRB/a9OgdGq3JC2bk7pCw744uBTSuNB8MY3fDpK
2LoDIZ6fxkhWGBQZA4P/xXP0VBxZ4iAxDf+ISTsJT+Bz0xABB7tnATQaI13wvcjemTLZaVifrAc3
BioTwtKzpTcQs/kr4rLyUx7eB/cZEMUe09UvFgSO5X5slhG2nj3HgQCJoEDBFHa53HG4Kilal5Ps
waeOOATjk/AnZ0QTSTJss7LQcRB8Culc4oenfwCVGb8p54TGh4qVYHrnCfgs4pABxFzYtJz/9xvT
4RqBxBUhaRToK4b14BSQeUBcrD0YdSQ3vuY6Ny1urfdSvzvS9XHhQE6/RG2AndZJ42MTSJ+DhRGR
8p/YPK3/3KlZTumRR5+jCnlgc25yfYj/qo+sB4bF8841Qzh0ipT3rtX3IjbL3CqYMb1lbUmvHbyl
+PvRjfhu/WokI42ORcZmalw4wIDeGfrHICkqo5kUJEDchKbBf3rtV1c+HH+gXl00GBftEN6DcEfQ
zYjhLonytXeopoqwI8yiQvyqTCxu3b63zDTtfaoGZanbrOVWv5IWw/azOqoYBN9SvUs4y3zDtylD
jsmAtQL7KTC70NHLFm/CN2Gc2E4sTRwYh27RwgIzqFDpfGkm0b1CTPWS124hzOxYv9+eBx126KWM
Q7QcgRsGK/pzENyifG1NsWyq0ticiQrzxDXDkOasM3ku91FcnwjpgjVW+iHp/TO/NUp/ztxIXAfr
4u9lsjk6wNwjHQQ1s4l4JtsKIpu/OZAf6vcCM2rcsFAFDFEEebrDfwes8JoSQD6Ps0sEipL7PpER
2uKKF34CuFgC7StOIN8dFKHwm97eroTJ0l/p2IyqlzbCvJD6ej7911AuvXS6WL/Y0V5wd+Cmhc1F
61gsDdUNah/w92yUTZERDTriw1YYoTpkn9PUmCBz0e34QE6XqPJrqdpV/XCdvUCtNCnhgmBB97gB
XMcKKVXBRv5VijiSleweLxNbz5WXTQHAv3OPc6LuVLAT7veL74QnE/FC0ESFagARFQPdCiMj84Jl
npz0csP5lEh+da6YvZaJAP/NqeWFKcBMvCRntAzi+sMc/geUeBHLCSLtVTKCxhXV5bg5gA7TN5bB
I8guCnsQAupW2siAocMMe7WtKNqHSfu+e+BO0NWAby5k+QFog+OpaqMZoBL+Mm/zlxHn45GNHcqf
viCefZYH5YtBihhbtvlkh8ozDqjflKwXV+Z1IjSeLL10bosHv3l0FofsPi25A1z/ZnXTp4TuJVSn
oQ2c9AwATGgfVipZFxJRIEF0BaQCXYdQDaSEqSscEoRT4lQDbI4c1SlsvSSUO2gg5tL/nShAQ22S
SocIWktGg8HL6BhQ4/VAvIuR/VDM79YX6a+vDy5WGsMQSaGaPhUvva0OI3L8yqFBTH/RmQrcLR73
43LTlYGQVvNc+U3xz3I3pD+lM5cyImQShpxhM5DX7WCKpGVuC9kMeQr/6YpkUxshSRRJtgKlaA/n
fgc+dQ3fsGW4R1Qg+IMM9AtyqBjYGB7+Wun0e+d7S3y3NCLBv4SPYRtneUGrCj2ZZTgPrEOXvj4Y
VULMCmyqEeAgPeEoMGk0t+pEa38HSeRV1UExVqlPAXGNv9Hnvj1HL4k/Rco1afsN6Bz4x9ftuoLx
g73f+paHlQgkmJJnbmBZIw4REySiftMnwQvhOrjfxuGCxP6s9q+ZxB3PmBirCx8gzzQARkX/PV54
oy/2nNP1buPolwWsb4iR25xVkQCa2mF9eUb6TP0aiCI6R5oxCibnLz14+K1udoKt/X8sw5frpAh3
56z3PzN7BWfLoal+JoPoTTORTxgJ5SIW/sZAvnPv5nrqIQKeOSQssuMthKrQK9/xvCQwesO2GP5W
gwlc5rbvjH6h+N4GY4sWpTYhje6s/tprIv4/o/Pd2Kn2Ef/yAZUhZWcx1I884qeJpaPDSZKkICCc
Aw2Fqq0msg/Zi0JC7fQnC/OALXy2mDovuXS187GzqADfCD3dL4yA3T+ll95VWN7D0SkT4QqyJown
4QHz+DCqlMJ+ht+/ikHMNVTyl+XUqHAJHQkB8il1EBUb54h6pQQXNm05/9Lq5PvMHn1/CgbkSwnC
jdbTf1SGvTqFXdzFANlya/QCAt0XixEkvVkjXhMPK8fc6dmDMgkG5lBDUvyInjqXlUy/1ZvNK0lK
m+4UmOGWyEKiTrmX7kG2I3Q0UoMaAXiJTIDD37Hec7hueLiXjpt1JW01Nts+V+/rWQcgRLriawh4
3fnQYcxBAGRfvXA/CCDhoksr8KtOCOma0ooykQbLfoqx0okqzA+caT9ALQumLI30fuCn6blGq44M
HZIHQw3KIwL72iODMgPf7Q0WgeIR0S75/uOsscyquG/1NCQglaR9THLxT1o60pNODMbnnFcS4Idl
TdG6QNw1M0kiJQF5T0M56TIBhpkhwodZwGHVx3g9BXE1VVyXYJSno3MvyKEdXOrnNX80KiK1SV50
jjq/Z+tTi53QUB2wNy9fFvv0BljIGIOdUuLhkAKx8zuT1AHI3gBnjfD3wFOL0K+0+vuxE+hQTNDs
PjqSclXRWDlOFBMIjJAHjzxkvu/l63BfYRK1ScieHKHJRw5puX9IKchBuDPwBZJ9FPJ4te4Hnoe4
uaweFQhc1LN+sHP+1hd2PpZMKZZ4cUbmQ02YTuu9Nb6ysV6Hn250hZ7BWiupQhA5UfHI0ktys1qn
upQfqCq1xTJzKZFJb5shCr+f87vPrck4++fTyR7xZDx9WfMC4sch8a7dMIKjUS1x6QyMG4rf0aOa
b2eS9XDYbQu7mmBVyiZ0YJTf3rCRtYXNxToDdjFwCyu1ng49N7WxN9FSoHuESJGKRSCpuc72HMvH
E6yWnsVo6c7q3a2xW2QW8+FvJbEi8TJnm0vm8+zZ5x++CqG6K8x0WM0HI9zQM+zK5lmza+UFiHkZ
K3/E2vkjEXZwBN4b+lsxW/A50DzN/Q9LS1Jrf1BaMbjgDvGofMaAttALTkNWj7vM1LK6Tbok6YJH
+N/qHbStXWSninbdr6hZfMLwOhfV7quROub9Rbb0Ay2HCholBQqv6RTb3O5MvGFozzwa+L/lN+GP
Sh+Sl9oCKO8YMDWh3FPdapv9Qiorc28k8mL2CpxWtn03qkxHQ8O3jeqEA3iLQAqPGD4SYi7KY+Uj
ELW1e3bLwuRK3jHIcM2fD5z7s8lIFMg6jY0fnVMYjAtTVOt6dCIXcibw5iZw3m1k1I+HQzLPNslz
4VINfEEax0B/GhIZIHPZkbgODbcfDcJ9CjwBh29U90fUhc+DWVD+F7FDMX9MEks/fKNKm7FoLWhL
YqeDtcLXnqOBXeOF3f85TQBQLO2B4ZHp7KfJNcV5mzkvzBKtcGsygHip0UeP1DWkzoTwDhHPqX+N
6Sh9RSuA54faC8YO84WDRQr65VUgKn0SJrdCb2UTqh49hpBB/zNeivzQqAS7jAeqTTfPI0eMH+fh
Mib12JIZKyWq1/RJBxhuKeOcyMmjEXrKLU2S52T0sOa4+uCRYQ+8lhnotFEmaHcLQYHyXVr0IAcG
Zm2XFVOBSP7j1a1+NPJedpkV2LD6csiBTVD7mQzPxYqriRA4hlFkJQL4xePT00PNkb8j1SY6NY9V
RexNiS7AJETvtOq9cx1RxsOzXLiWzF5MEe6Uxwryihn8tVilFet5SegYB7sCCsfEWrOA47FksXJO
jdn7w1qgWADBLJvua66fvvMZWqF405RW4ScleiH8F04lj2FWdmYfIUsEtIktei74iqtVVmSd7yto
tjjAYGjpf+BXa4Hr3w00jvgWWaaYBBvvnGRO7LjQs+tAr8pRQ4t23FqOob7CT49sJAIpI6Oj28v6
eC+Im9HcIAubjl6NZRvBjCgnIpRpmIwJxOFlCz92w5L1DM4NA95bn06dSGE4A6fne0kkaxEunAo4
k8pdO7hv/OEj9fX2o2HYajV3eKH3ven/BntkLXK6OShXtSGRZkNUDBa+KRVC6eu+VVN34zwegqjh
s+vmMmmUd86c3RlkLFwQ49AKqCax7WKYtOCdJ+biWgEXlVy+6Kv04oAJGe+KBEQ0Nf3qedkofJZM
sHzFdX9ruLahRBsI8Gc7YiB3p8h/zbc0oaSSKE4KB3A5+VUITZ3AT7SumnzQtiKbKgDCx+4DZtNh
suZFZZgY8RbdOycXHqzeeUkqHlMFeoeGvHRuxPYDuTD8pWrqI6F+ZfJUogL5LzS0dZSRrmTkHYOj
8B4tscg1NKINhPlV7WWMAGXSXpTEa5WPRAy2vMTwMNZbV8ekTgvbggY/2D40qWER7h9EENN6iGqK
7gsYNzJWDVVL1Qhy6E9Md7Nyo66paSiA3gpPpOCgAzVuBKJeEGyiHbvVl6ptgyOZdh5HIh/A3XA3
GSWslmfxdmLRYYqeQrTXd842UCSaUFcZpTfSOWM2Ho4NkdZtbx0WPx4ZJg6pXd7aIDOkfdGHR5VJ
eHpULXOd+0jDc5VJXqPiF2TQGal85BC7FjEARwd4Vc7HdUkJq8QE2JBPnLOcwidx0K3w/MZtCQfE
e72GqzqSJfp+ChqqGGkGv+LKvN1KZ16dY9wAA7iYutXx6hBJEPU5I5/GYtks6H9b18V/2CT6Nxpt
gzATKpXBnD2rA7akf5P4YLSAqxzhNdvoOPPOylTKbRHoN54kV2K9sSgKguw5eIILjrmPQNoIsI5p
FSlGhYH8WWzV4HLu3hyWxPSMH+FZekJNKqaL64uGYb6wl7u9mtkpDJP8Cqp4hkxCpVqLwWEYJ7L/
E36Ynx48PqTjf7H1K1Izx0YPrBU/XHZMS2/SRw/AT2ZwqzIaskcS/AM/ibmFx7Yl2jaJLq2cYXUx
thyhoebjZ7k+w3yYUKI5Qrl3SnlWZ6X4PS7xbcL8c9VaeGU6JkaNcKPHEB5yWJl8avDXk479RGQ3
X5nJbb7VUo9mHXiXxsQ347q5shfF64rYOvGemv8+4uIUTCzsfwXTNgIuvjqODWzmjLwKycL8Rse8
VSsu+e3qY4FuYiHQpjKBnqXMNbBMiYTTq7dXUopAjbC4kAtritzdEbIG+mKG/xdrXCrjR43EQnev
yeaeDATtJ49weRKZK+aXPZqQyn/T/atzINBG3muDSXnVcmc/as3vaXFcp9FbHfNZOruWTQhLnLcx
6f9TGRxLog19YPHetDtcVaLK/eofqPggSf5KAcULMoiZEOo471jASIxX5Nf4V0z4af8QxCSc1WKs
vBiwJ02gKMB6Bm6XHtujtOHyJveVbmaPIz6Ah5mEkRzykRtkYyiUC6yRrrjDdaeUeXHtyaQKE5re
sOIPDhUc5Jdzru/LqaFCl2aMdBUUDLJWDWVY+xd9Fo3LcF9Z0EIe3tQsWgE6u0kp7SOuxDJ2M5Sj
D85LMyvaExmzpx/sVJ4b3qS81sMrYBz9CRYBY7HiI6rNtr6XAIn9FlUBs4XvuBLttLL7zThD7WFw
e2ncQvozJi/X45eT8XXze9TgKPCRKwHek0B9jmaPW4Q2qLnL4VS+hudV6Yq4f6QvJsgVT//vUGjo
WQlGtsfpUmToOLVKhLBsPPYbzqx0frgK2Ced9UrV9FOH6c2S5AT4vMVrd9D2pNTxEZkGLQcYYVXL
F9D2uBOjSM37DW8hlX1FAHPqlf74liyDs6i91R9yYusPKSE45Wkz+OZu9h3t+5AEjIhqesLgGcqZ
9EkFYIa48Y55CpGJipGIRYwTTixFngyE3OUC+GaUrOSj+7rs23nyuResk9e24X/sDGtLKtX93slt
O57x/6F1Xg3jJEjTBG6sBktkmErurN+kh+SKW1+UsunyPpsS65R5VVBabNIEM9tDhjvN/eLCb6Ki
U7dbwVXOy7R8DeZG1l9DVZ7C4menhmYbCDDQ22fV92TscTs+/viDk87Tczu4P7ucGd3dT5CXTBGM
olRl4okCpi6vyCIawhG9f1H7J3mIDE6DMmONfHD/N9vMK8tkkXq/SuQ6CrZg1PW9qLpwY27Xd+g+
w8zz/cBjhaRrAZ1Z9t1MITOAfkGFf3qGXrMXfwiapgkhNp7rBT82GYrK3pjQ3F7IatKMtw3s2IEw
1/SUQ2p5h9yBsJF5c+ZGWXI38pFzNd8vOAigvd7L5nLyOIOGnWmrOlcr5mDscmdDXzGHjEGcfgRA
iFmi1BpquKr3nbykcYsAq6AT8cksX4R+TaVl3NQAJtwp/ijyZAvLJlbRNP/V21j3LPQv8949boXd
/1Gb1bdi+YH5/BeioY0VAfzRHWGyHZlFhY19Ogogez0kSuqneFtpBcFZABrNX1PQILXglBBxmy/6
j1sKnZeK4ddmZWH6l/FcS4odVl5WYmT6ry1WHLMFDtVGNQyjm8Lo1A/JAzTTJ4DueZLFiZSGrZ3Q
8hm2I/e+LaUyycBo67KCfo6LmxVBmb3SSgQka4KH4W0dZw9iuV55N422z6F8Q8OtthNCiNj7VeBa
PWA23cEV5nrTm8r/ah/yO5kb92tM6fAIlcroqwfGvZYUmEtSF8PLO4NmaQU9PknCQTzyX/YpC/tz
CYGN3DeoYcDM5RFi4CmDNzclVcNm2C1kbcLChBno7gIntz7lGWGekpNBfkrnWXwVGu2JwUhcpJMu
7e0/4Saufp+y63XmacHU42eSHBfkQXDps78KSUjZROJ4pivmB6kEtLyVi50fY8PSM93VtOvJRShx
m7UuTcSQ+qcQbQ121duodOvfGtG9KzBg+n23vAQX/z8O5UJoAL276YLL/NkT02T2DDC7tejw3yO9
/DA1zpc45ZKZVMmirVSKwq0eYWBS2mBcJv5wWEAK50uOifTqKkYPYeDrSJBKmUBrixVPFdssV3OV
moc8uxHjpvXWBjNIOuLujB+XRdQkPsOYT3wdj1zTkDm97OeTDePpnhMlKGIOWT/xNJ3W2jp4IDAv
e2y6D+ekkpLy/mMaBYgf5m+ajXwL85agHpi1at1FrWd0yXqkZElhfF2gAzoVtWIiOeH8EKRodBw7
U0kFFg85C0rULLTEzX/t964GmpHMio1ATQfIQXLfnAkhQE4WNko3uOsFKl2FJxcJWmzFupNBUtOk
kw7IUcb95yLhcVHXHQA9Ib5V78jXYct0f7a9a7AVFlwK//fCGhVFVtuxoh/76xtOPq0viSPthRTC
hj2DN1jLp6Vwpt9BHwtWAYk/QZTSgR7tQyExQ/qyHgvbrvzP3c7ATxOWVryCH0ELgKgQbFsBYDes
Z5rCw2L1goAotEEbSwPKeslTmq8uUwNM8UURDcN28dObzrlmGFEQdatYmhhtuhfhc9yy+horPjJc
Lum9x1duMl1nJMyVzpmdE3nQXm15WAsO83pVxPr4K4dr6rNHdjvKKkJXqKHpKoNRII+p6yMOa1OW
XDO3/gaKu/2HJLvYqEDAiwnqQt7Wj+SZIXg9R90G9FOlFt4xNXuyZgkdwvBqDLFmAjq9EpWE5bVt
XBIBTXMjN+SaYPSq6iYj8DAysuyO2RNMWwsb7KyMH5IlJ3HenOCgvtxR73JYSgjO2G1SxhX8FxjQ
H7AXdO2WZtAw0EaHHbSq+91JgfqYsBCGfb/gm+rUa+3Zq+y7Y9CrlrqIF0HGd4UhpJqfAM8P0JRW
9VkjW0G1tBTmTRaNYxljCPcF+Mhl9K+/WdulnkCN26xpONeGscMqXQAzgmlBVXTVj5en7Qg7ypfA
HkmqFBbtheyg3GcZk/0oKV1gVBwvF4yMIkYul6sQSXDW5cpuZi0XCzhsCcSg8t3KIgDaTgsl1I8H
wAKJS+MD/6fVW79MN2+HnHRREFowMNow8COBUBHA6uq03ZzJzFCFPivPKc+MyeDaP70p4ExSwD2X
iCoq/mrHCsR9SxZwC6O0xXDvgOqcZF6L5piqFArn7krr8XMDLO4lDugLREe5MVEd5v0jEui2RXcw
5vqliBMBiDJD5+PGJ+4AMA2yMVDzohmcco37eMwn02i1yiBVeVtuFS6XiWkfFj22Lwm5VI0Slgz+
TtHYKkQwJucfGIo0b/YBdTy6piWwt3FlkCMs91tlpkqlzAKWkrG9lZs/A1yAmTv936kmMLfF19sz
XOdIPA1PzkHOuwFH8MQKnDjVsuJkJ8NA1nYUNpUqhf8sI3YfTOq0op/sO/h0AqB+oYtGH292airo
ffbCO+/jh/TYv3jhNo5ravsh8YY6CS9/jc6OzqxxSi9VYECSeJD9lzgi9LCTzOv0RlrZBc/JK2lz
phEs9uJMHGeDloL3Q98/5FxweK+fAQOnf66UMXwjAxFBJs4LUo9Et0SBq8Prm0yvnALHmCjpbbO0
lKL1LQg8N5JYnoiOtrUdkxFMzG4RbPX8Nz+rcsDYAEuuUW5q6CheUXFwmcztE4SBl2YbHqBa5rLU
tOaw8wRkXbi5cMJe94JFeBsboyYzNHEVsP80Rzctkyr784VCHUOCQwAeDzJSkvDxpeGdGGY66w54
1kF6s7I2a2Nej4LgDuqTPw39y1HVvoya6F2DaVhJjjczZPY9VU0J9iTDnTtio4/NjzcxAMCMb0vI
tbfSziK+0D9XGH22snmMA7DJb5mzfkKgkCsUPU4wSuZ6egKJBrzbctBSvY/Qy1J+ll23BTQYGoIq
wHnzWdw7bgxdmzJ+hYIza/Xf2UVNV7pQLJXLao2ZwDqLKf6rQZNlOobOIdNd90j1pMU0lfSC0ihy
w+ugjIQRLejdSwjYcqHuKcOzbS30CciOyRtNKzN5199e0ywYaw1a+NKdTjeNV4fKVu6ngmCp4jdQ
q1t7e2/vwfM88mjf8PXzkacfVYQMPbuI/JRRGBGaSGrE2lj9pFKvwmiMi4B5ytdGoD4PQt9f+uR1
YjkZTDVJlhJSO1AjzuB8HCmAvbgVu1EM6Kp4wNDz4EOPIARV7hvHtf+4+VwGW2QihfpCsBlaB1vx
SZTaz6IEJJxO/fk4EGvtdfP/WaL/BATd9W8ZytnnC8hGdTmlcHtW2dJldc9B26+p2YJ02kbFRrDC
etKoyXtv9f7H2Ov0NCLfAS95rJmFbse0Jj9l9cxo9rOXMIWMvJ9F7ySV3rcYOHEPyDU7LxhSE0kO
V5+wZgYijTSNVP1x1pZI8BC9yjVLW/B+NxIvXFKQznl/EoM/YljuHUv1Ehe0syIaiuGXdQRdfRUU
53PwPHKUgc+SgmSQOSbMx0p4wL3XN14LDhBwvgISb1oApvzgB56SW8P6W8r8C+8uu8FpaJ9IQ4TY
89LTDNKg7E2+3b+B7E3aWHXsnrxjMg18QKIXu93I7WIT7eawd9z6Vdyf6V6O4SK7x00EYpJlEPuz
Da2N00OWQIh0RombucCAWqpgp+/cnK6s3X+3AyQRfKoWjdW3CurfR2mXGJdiWzM223KhOXMulAeF
bXqgvK6KKnUdQfIwy9v7CCVXr4RDzZOuFNBdHHQlPlbS79vd6XnunKzQ8dexfWwDvOfzMjT9twVm
6VR1kEhtyCW9ETfAQDO+0csY2vUyEphLMXWdO3LHU2PwmYnVOAJ75YT2YmnDUIiSGgBXUMFVZgN6
ZFLk7n63/qfZlA8UxqOmiQnON3LFFKFLQjEElewa2GnavENsi1ercudvtLaE9k3XYutJSvY7zOVQ
e0XmerNWJBHOg7HeEzK0rJWDcq1gCsQdBlS+Y7BtQ0ccTFfhGBPFz21GLnAF8i1Bx4gwD2GBjSSg
67Nq6Krm8twXCs89RMFKN8gVZjz59YzGKej2UTOMF0aPxJkcB/5ULsFjQsQpPklr1s/AIXrypnnX
nKA10CW+llrE/F2q/J3duq40NfQqsc4gMJDzTcWesq2Gt2I9jMzLoKYCuQrw7OZWi/M3OcMnS6xh
W9yXOIbjSR/zxLM1TQsMGQV9f7UVld/gqF3/G2CHaPu7JJSQ3PiQfSQt9gixYG5HLAs5SUA+9+DO
yPFqyMlVb4dgXC5KaVQ5ZdLWxmfk/0+vtHH5MAg3Zuuq6dJwUSoJExhiJXwmEYguXb5JSE6FnwGN
7+G94DkvBRkjgZP1zumgw45mUH36xpFFjiJYKEz9WhgDBdixgSA737o78qKqRvmzmPkQX5DOfUVc
RTYyQ3RXcnIMQNX3UBr/afgOSb0QrGl85eElboCD8iNchhk/Oyg3R3FULpQzX+6Qt4DBglpITt/q
0WBH+OTv1KyuaA39JmPdPEbBzisT9QpX5NF9oAGoWlfWyZcrZ2e/DU+Yt3tPqHN1b2E5wBueKDb6
SWC5gfAaXHEim/desgBjFhRvMJTUbt+RFMbsmz0jehwoUL2g/w0uNLXfoOyPAARJADlJJzhmfTfj
eaO1IyotOBWdQS3RbTUbPnqOvbC/jslcXjFB7acU1EpJA6vHi8gOiQ46M/VymcsKhgKtLNZydgnL
aZJ1fqOHQx6NVuYTw0heejt0lahRzj1WzjeorYhDLBvorhBKSeZbrWM43FaNvT8yJeBduDLQB/2O
4nGCAXBWbUkGgK5or2Z12GDNPUL/z6IpHxA5bE2vk3n2psaahLrHMDyPmdaOqHHf6GpBEE1ptRKn
f+xh4u0WI9JRUYLuIkYee6aXzdVhsSv7wf1u0smGiV01KaxB7W3U8MLwRlKzkvfzO+Cz+Qw5QMsk
opyfywasIPfFt/5YkeaB+vWY3EmbG0TgSCwjgMghP6lNw5HMqbFrN9e87ijcYUQMzNyoxWK8/4Jj
UvQoOJZ6Et3hPqY65eV8l7J2qb7x/GuTFW+wzXkKVdOMXmU59td5xt/kzQhey6tB5Gyh/6OpJ5+I
JcUGOK354kH0hoFSnWlB9Ov/2IqAQ4bAR/w793MLEQzCMp8VnfTkz/6kokeU8XJvKSmVowuvfFg5
Q8s2qsNaXwIc5RJ0MV2WlSHpSLZLcwWpRpBRW+NY4cMt+VIW6IGQxIY9ij0UCbbJ80ib5KGQUCFG
FvoLkRNqTX2xlPD80r6sI95qJQ24jftkTwNDekeQ+DBuGslUN1JrkYW3j8QnuQHzeeDBKxu0q4kX
m2/M2j13kTby7Y3LFa5UXNab8LJM83aiIuD8rcuWzveKkBR4dqJorxhCumYB4h5SkBkuy4FgdM9i
hU7QANCt57yUcKB47d8dGByA/4mUmOyZfksKsn916KVDGeagcVsoqv/mHFzxfncptTTPsSKN4WyP
JpIQECor+41h+VRMJG6310/lFz4HSTxbWCefq1fIuNwrGcPjFiwT4gOUj/ONTXA1PPqMAkc9G3L4
7BHJrQFvnm6KPoV6pkEZf/rM5hCM8jH9vBUP/pSrTaTzNeqxhv+QFKW5y3TrMw0w/YAQJIJ+2LKm
Hs4z0WVBqApELJCBNTeAijGUcyF/buaztRGPhwW9edQ4teE99CPSj/gOBH3ShkjNsKR4GfS7FOHz
WcEmRi5ArioswgN08zuuWkeDqlZ3sgACJ4r9tsogapkJNaGrTKiDnz/LSqs1ofrPVSB8PBTH5ksA
SL48idPvzCn8cBnivoOtcLZ0QuXFES+OpLlMSLgRE2aXnNYMGOfqNJV07jn8nYdo+0Mg10MXy9/B
qvSEEnzYOmZoacHtoNkJ8OCOHTFwEpCW1tRdC9krRoGsta/eQpzfSGW2xcm5gyVRpPVYe/rCz/rV
HvB5M/WTnGWl88P7MoKNDqvWx+4g1SpsdfEB9ovYdfDx8cVRu8VA2dOVvVC1JgFHm+wcteLuI2RV
urk0KxCFGo/JmVa9q3uZM/fxObJlkh/8ao02xsD7uhw6KYlD7YRHiNqVKpBIBUankv2gXfaGwmJU
S5mJa2MEZcVds/xY837yWgsojFDnQYPbN5SPji5/y3XLS2Y/+u0vmNfMKWG/8sexDAZt4AQzI4gw
ypvD04OqSQsXF3ELm5bapJkeEB2YXjIvzsaU/Zix3PH1f/7R+by+T4vHJqpEJXAULNyL9KYGj4tr
UEvdJ4ac13owhDXm0xFOP3otNIQO5H0fSRquYoUvnRGF5De1jvtbZ4w3Obv28WBTCB3TA81BGjQE
D4KU6Xmtydyw1jQ5rgVR4jArxucJC9WsswTKTm7MGlZOsuvbmGqU07peUmMEy35aPdPHk+hLq2q3
94Ei2SkiJ1G4ZBbWUqTmlIrj384PPPz2kCAW5f5SW+e3A/ikm0RVHoTyLJF+6MejJqyNa7DTAGzz
QVftXEyIWGhVsvXK53pPsfBLIp2k1OW8hGG1SxcoBqqa3UdkH7iRBN0t+OJTEeHhsXw2XAvBrhrt
GUEeZ7wRFlUiAqmgx4OYnK1fYMUl/fG+cJzJSCsljHJK/SvfeZxZUEKxrzdgyFWW2OEAFR69hmVr
/I9mu79xUFewpHif0QQ8uSy/jhaWsmqVupwS9vzbZ5W4hjtrfevcYZ1+aatk42AbVT8YI0vwhvfT
mSxD32KLNGOxKwtInNjijPsWUDJl6BNEbZoRtvllKADN+VGgQU8hhmeNhhP7qsv1rcSDKmHRYDpL
wXr8la5OmTROd0TkohCouzVnBW+A9gJw3+JUjsoo6uuSt5XqHUD0uJwGeKv9O9qs8McHONS6eezg
aqqxujUoSRLmdjTjyuKjyzBOFUm3mkDCDS2cdtBz6qiB7bme13VuT0/fIuH3J0YDlD3WTTYU6JbJ
Nm5Q9aJaAwmGYSxdYKyBzLuC8P749N6uulIaG1Dpzo+ZDaS+iQEkW49Hech/gAP2RhxalJYwg9MY
oXJueS/Lb1JOLp7Rc3yFuP3VNE/D8VC98wH97jhS/wc875Jf0eE2AJdX98PfIqMgnrWAhxRx0WC3
DsVqcQd9ZeFFxDqihfskjR+O1ZAot/y9JoulZqiZ8oFEprZ+j4hoTzlRI7rBc1SFcyVVAjj2v6Nw
DehwMK8ePz2IE1KIkNz7T5El6ybhv2pVCNm3Jj4+XX4RZTtHYiiR3zEzb/OWiRUZB8qJRaryYvFL
/GCJBL/AE5TUZlkenD6o7dleHeb6OmLMMW1jiV5vuG7ZeGufNuG/lIFeFivqicRn2/Icv1qovleo
GNZGPX+FqN4sWeOPoc2k4eyIsxEL87MZho1fFiAM3z9QQEedoby2rZKomUvQj31/zbKm6E60L62H
lBV/iN14e/avMJ52ViNxl5oEjhYpC9Y9N1WhV7of0cE1E0zFAYtkaEb1CSCrK5kY167zFiTrCN3Y
ys2qmkD+ywKeEvBXPDcrGSPzTUFiWZph2sNQtfyaVwd5mPk/JLI9qicjGgguIdHuWm+SaUk3C1wg
NwdGODxucxaReOLBVhkdtHq2G0pYKf3qscIq9qiw9YLWOO42OHzG53n4D3toZLtv6ktwNEzamVDV
hGWRg3xypJTlxFh3hM83eIBWy0L91E8+vyUJFWqe2lUL9WIGLawv0gy/Vs+8ScUaODFWTE+R6+K3
QvUSk1S1Ofh3mVJj8xOTkV9S/14DTgF5+w0gLwgVLjBmM9JAhG5wSmAL7hBT5/g9UfbqXXVSGCmP
Ow/7I1Vu03jSm8+DsUOkMutWA11K3Nv16Ncay2N7Es/3xi7wu2gK59m/vgJN4N5EJlqOytFdmKVG
vCr58+/wIEq3UaET0P7m2t9DXCA8FK0qWeuGtFoN0eY5Hov4IzgqoL9QBdc0cfH6XpD1liudZXAa
jGKx0rjvFalmIw6nr4ovz67l+J5XncBOtybLmeVzjXZ+nK4pl+DaiJsgWSFgW/wPJ6HmmGsYCOg9
h65nyS10ry6nZicHXfdWjJ2zj3iK5+3KTDktgpnNY4nQQHmwfHVS3+t8H5Ynti9mjt7WF1i/hfJ5
QENY3AAD+nFWs7pMB02Hofqujtk2Gteg13eQQD1/x+jpgpAeaz0ZBuyy7FJW1aPi15Eo4XOp2AlF
7g0uf6dg5oJ2eWoueUiElLUfZRRxL0qgK0BDV9pVm3dkjxnYk0zX/rsnv1NrdANAihvMpIBoOIi0
c+mKLlGY3wGx4Dtr3JatSETVtXZWzXD3/16wUbOSyjNgPN7t9cjJi6jcEJWzmbw8orgnBX+PC92f
QL0clmw3b09C/vjkbwAwWvNtWAw4EzoryEHaOPs8TJGES4X/xlGfvyQ5+v2YImB7UtcGcP5gZDDq
GBWQDFVKLrBOb6jdLMxTntDPETmaTGSeDgXF27rRbfxj1X7SViL/8z5aA1pH1VRllw8TkbVq8Q/T
yulOwtH/xS9yRnvhPciYyXxDKw7TUNC8pIPL/cD1PNSvE59KWPMjF8iAVqehz9dMM8SWKZIf1eJV
9O76oepfX4N6j/T5hMENKsAbpqbi1kzeczjb7Sl/LiZs1wnshJi4Z48ISvg/4UZbqH7g8xTIGs//
OOIur/I+d5cbwUtlP41gzmbiP7zPxlYwgKeSbhcFElzebjY7eaj9D7k1/DaBp8VbVeinCaFU+2hS
kZi87IYOQ1ljWnTiA60o4lyWLeCOCYjwF3WeuesSN4ePl5FJcneSQQncfEB6kuOfsVez7eNCbo19
6T5Ah91P7KL7Q99Wje76iqmaj8H8x6qIrR1wxs59S5hWhk4uRplHa7FqDasLMShHROEJ6B9f49zn
2fxKKejsALizP869+yzns8t36IwqG//33B3TMPUjYl5LfHBBeeNhgyHZQwiRUR+DOxTNNF8pRj5X
BQBog3REeF6Gi5A9fMCYiSs7uMRm50uGUnGICi+q7PEdGgYX1+Dc7UCnAWTyEyFgMy1dy7BjKVh7
j3Nh5rO8O6f69hQZqXkufPyben4r1P6mS+cEPKtLk0xwLttFKh61VhmOsqFppOSUjO8+DKc9aqu0
yt8fCmUkORrrPXYKR+zgn5/pApeYkZyHHd1QvBxYis7D5GNWavnXuAYwZFQWIjKS1z5kOi6lKfJX
MIGcfD4qmKJ0VLjSU+yY4iPKSWYosAS7OZEpRlQT0WRCmXNGZ1kvdEqHtydPOEEXY+IXCPzVBB9w
6y83L+O9QwCpRMswPMuw6CER6IsqlPn0j5LjdSuGcflQob2oUlOgPkEIKpkYctOA++zEg02gCHZE
6w7T29rzpUKaqH6mw6sSZ/FhNbUqsC/poppCknAliMCbOmx598C965s6MLc0vajnNaxeuujTvpFE
XjD2IsqxNwvKAPzys02O4s1YHYIimHxiENpOErxHNm3b3fh2z2OY4tG6tJSo6PfETpgfpbSuIB9P
XarFsI5Y2W6I+QLZRNXqgUzcEmldYM0Hfps3QPeh71VTo5g/Gkj6IE0h5j8OTdFtIM1ImTq6ELqV
sRZ/nwxPgUReeY8ZhRdpw4DeV7H6+aayDrlO1KiLF3aNt+xu6Qx62AjLax9krZ3tVMZzMeqFPIfo
kPR7HeN1dQHjlQPyEZPsNcilGuvmdGUlaCejoKdJSgZEUFXWN6Gg6S8AoocOAPm8UwA1s/yl9r6c
hZh6v6WxazEROhdiMnDVBqk9iOKdg4jjDeGFj/UcBSyovPUhlF6nFbzEEK5CFO0EP/Mqc/xub/J6
DxuKuOkjJHrki9VTeGnT25a3gS6BRWQjjMgYVWZZJB39dMF+h36rLnVpQNPDl4v1SAqeaseiekE0
D4V4yAqrzPsjW7wA8vrE3xayTWhjac7FgnAz12qOehwYoG67IXXmlp9pwN5GKf9oBsfCagFFnrSt
DM5tWqNnO3TiNUvM0DBzh1Y1YOrOmQgBsFW+SaiIxgPL8O+WvxQbTcsFp8OdE8okqXQg4jdGvF7A
rJ1IYgMOC5vnOXP0YzOIJXUe5i6G23ovZzALLP8vWVlPWOwt6JigOs90N7U5vx52GliMstfZJ44J
EEKE7C+YF14pW3TUvID52sGao4kYZ1IyDwjYXCNP3jKOQ7T4NcQV++tHrOeU0KWPpyFwN+ZZN3E3
Y9iS5QIqeJrPY5EqB3ELCJ7Ps3KFJ6QZyT6Pc7Hh6Jzq/HD3KNCsmQvNelAtacf14YfDhRC/JvaC
U5CpE7oEQU4meqR8z9yTxM5niDLSgGW4Z04GziyKvAH0tM8Z6oLy46qryXpeux/gDCfjY2ggIN/e
VTe78XVF17xNlEuZ3IFC+tTbTNTqkQErbcPt8AXuB91OsrUGaPHxhR/PiAnqA+Et7GQJi9S+lQ5Z
B2ryT91eHN7gvD7Q8RG8BJccG4yM9ze2Ax3eO/gETMHiA1nr8kK79wSlKK0VqoLZ9y9vlL5aGZ0g
gMAUY+rT07AdvfnN1rqUgp2q4++UwbU+s47jOCtEgLKqXDNy+tBmdHwBh1+F+98qjs5Yu+9AHKMI
BRtNIcJ5oSmc2s9AidMsY35hEAS71thXGLZUip6l1mIl7j7AjxPNiSSQqBmAqdTrmSzbpbeTahS+
cA/6Rd5rjCsadz92UPWZGcv2+Q5EHRy+Qd8qyyUvLb+QwK1xoPFi2ALA79HqOoNnaHW4XUCjr1KD
s91mgxnz+XKwK9bbma9/YMd0FfebpbsU6g5vFfLWjqGvzsJ/ZjZ8ARbeiEIs3LSJ+FcXQLlNYVH4
6H49db44e21Q0PbV2nt1uTXcRi0cGOfd+ENUqKH0J7X1Xgz5GZiostxgFgF68Vwj6xk+GL9ZMyHa
PfGL5v9+MU1p6zxbm1f24YOuP8z5B84n99ar1uJhZesndiigVjWlUuFCzp8b9LnOHKqwYgqKFtSY
W/dh184gYgQTPHL2/Cs8WXC7BvSgG/xcLBAeJDJMOmjpytX7vFk15k6xBMTGPYj/IXKYwF+mT8Nn
Qa932W5YanuYs2PjhBZx6rzK1oHGG0DwOg+xKx6wI5G+XT5dyfY3Si2IhtxrbSzW5liuXWDjtsTw
aEHXCP8pEqu7w3I6Ny2+y8Le1eTYbt/jzekfs9KZU6OGO2QM/AHfCKyN+Fe0fRDYAAxKiAOcg6hE
p3vDdHUyJ/clrnEKeG4haDsMSqAM+CPUjLtPfuhdAAzbo2O4BOSa7AET8/ZkHDxrEA/XN3ekYyqQ
SiYmaFjxFl06XppMxyYqPfqi9VCgCznMw1yf05KZoacbUKMSkkgz/WlEctGbU334Buxkb/OkzOSX
ayc/99UEQWvgwLNLMvaL+l/eVFDuOi6otdfJ7ruoGPM16cUl69piECT/p03BZzZUKucaSrnJD8gd
4tJBRra9MPTnLKG/KOAJ5jTjYLyCHvqFGXmL545G9SjUWilkvZHUF/zEc4D0cobqGN1AQncIXf09
tuL9XiyTrO+45IqMj30TSUtjkSRUWY1iys+wFDUed/RTm4oYwZBvnYubC5BOgQYxa+2+wTuVSM++
g829Vu7p+ILHzdAtu3pel2KGJkcDtV42tWnoQu8fbmVznpfCZTxfyAFT2IVXHSckstc/61NV8D+U
Tz43kwHSR/qTq731JzhPgRqnB1B4F94MXWkimQsGkpMQweE5aNH2urRHnQgbuukyBJlmFdFamyya
UdHAzi3xbZCUe+d0o+Qvw5auTZKHu+1NREw44fixgA9Ep+OCBO8gHAmCzhqhaqhOimhBYTWqvuT7
HjqTEAIfB3+1CkBVMovsMqLDCYvgn2kEZWh1SdLHg6i6dUknPISfwQSuKpFsJ52O9JyrDE6D1oNg
WkYTfg5sTliW5dkr7Pdz9fAWfrMTpIBMPCgK3G/ta6rczYdKPgeyazE40v3W7DGucjVnv4UdATUb
3eu0CjwZ5VTpgvOwu9LkjyLsyXobxVU7VIpBHpuOJY+75QXPOqdLwDh1iEtUfYMoty/lUwGn4ZqY
GDQG98HNUwxh5jq8qhYIAPqfFGrP8YsauGRlS0mVUVMSZhXtmfpvsM3R19VHQ76BnlTWqAl4wEFR
7YFI6P0jt8lC5y4nBmMZarqFKnR7YouvPpWPBi0JKuGd/76Vag1mESmsSa5dQNRlTFmWRvew3doj
gKztrrqYXMkuNnRkdRweihHZvmR8WFai6rXu5kl3tlvlz/TBE2COUXa4D3403HGlSxKMhYxg4heU
qb9R5DuXV+oxCjEadbUf0bmZSJCNwDW3a4SY6OdtF46JSkYNcUOUEpyJ+m2v7sNGzTzLWD+cuWnt
7Mww9y3x2TX6Maf7SNMBsBLydDeHQ5uEMLfECRMouvhawMqpy1FOe3d1EYgneR5w2HulTQAjkSIw
ENr71L5+heHgSmEa1XENOL2ZufBPsX2moUgmRkehd/tF0TLZWAc16YZZGFnbl6byYnx/IPS2lEh8
d/gjNtV8AcaKFAaDyW5+FUL76h0TZ6er1VyRDTBHcQXZvm5dB0V6fLtgaq9GyR10DUDEFr4uIubo
qlpFYpUgGDu2t7WQtVKVkfcL20cTnhtVfxQ9N5T84+0G1ZVrUVmi8wdhh+hE/tn+m/+l22ZIlwRa
Yc5OzASTd2ORMg6RLmAhXacGQtnloD1QQjZkp22VcKHpUl5rLgXdHo+hcxCLH1tIRW2GjpwJnju+
rqvaKa9yCzM20bUspgtjQR6eq8BAzpUAAMV1SBPrif5bX267MgCt5nA+J8x+a5yshsR47JT7Iesb
7wNCLwADaXivz7P6DmC1qUzLf4QVthnQJo4XvmwyjPCvL417FMECthyjadXjWva3/Vbj8YmoRxWp
ZoeoAlrZQKLqE2I6WdQrKw1FEu/TSWi9qQutpooxW9BO/muaLztexQVQMsflqxbq0BMjnAExYSTg
V7rTUivt7a1pWtxE6ldjUtT/NXWTnmOL4/oMm5h2UQECROVTOIV3xdPRj0TzGrzyD/x5L/O+5sC3
WhsY0Vob2zUc8oDQ9yrg2pNPbvNUzZqDYCzwUICy2G8H3k98J+SoTIwk4yNKGHBIVRM4Qpav0S9t
kIXYM1H9QgIAtFC1AbU3yzQFcYVs1DIrb2denx33GUwYUh9UgyvjEaKUl6aZAyrFwJRJHv45mrOX
1bnuD0wzJKmb9/YNt7Q7kHMDGKaGXSSgRCGfqemLSgCN4PUA4u6HxwYdCDCpHGbykm56NOJd7NBx
hbKagZHupo8k6vSKoz2QAoAzJ1yU8vJH8XSEDynuyIq7YFWDdxo2XLOVtIlSiY3TaQ1/oqKmIgC/
ktgWR8wvFJMUGO2ZUf1QgfUehZjVKr3l0M6hFYSQ8fGjkbY9gBcEwDNceLtB5t8/yArBPHR+E9Qp
VAjcaQ2LgODlvIYeD51+0ggeVNhcj/hwEiECCbNXIhVv0VXh86pfR4H54Bwa+A2l3NM6fb/iJlVC
3+lwJpi0ojywfKWYthysayqpcp9Vj9xGPIEXSKAQllxmk1Xwcj2roj3HSALy9ZUfcEvGmX4Ypo/z
ytwrm4K5CMdddZ3nXtxO9C2u8+YTsymEUKXGHBYSX//WRJp3qr6mQWZrj9r1p6j9Mxgz3xjrC85B
jqXiMwlVzm0oJHKiFrrQmZ/zd6+eINNYxYIaPnPw8GdRRlEuJlknIUbr/+DWW6XwL6PpAAtJxOKq
ocja5yVcbDps+h1Mw6SqDKp2uk9KTxs9n6EcCrBM15Z8NsWnFqmRpVquHiklotNnwaznGg/txFjI
LLo51ITEA5sFKtujjHE0jIWmjnXE0lQJ7tF6wjcP5CqyHW9IJqP+WUUsYdk5dsikXsnmC8qx62zt
PVR4laDJMZsBhTilkelHjfgdOUVmY7bwFvpt+qiEPJyPzQ1/1RwR+BYaFvo21Jn98oqwXnoxDw+r
N59/fHXw8Wy7jHScXsG+KAZAiFVBYcNNaYyj/FmA2Ez91bQ0pe8bo5PONFiANV6g0KcBEq8N/lV2
Gw3d1Uhz4NnI4NZGXXU7xVxWUFfGwiHtDEbFDtkP/Nyp82ZvWHwmjrHFes/y9E6ogQfRARZDwryW
rSfsFdLjxSq0WG5q2oH5egBokax4s3UphHlXKI34QSPqne7V4jIXPyls8mom0n+E0Ma9L39uHwff
T0iusCat3W6uxxLy9KUsL3JVj0LUeDGNb8tCywbUwWeTE7rs3eTuZBvLwp9LgWHV/9erLinjkIhL
FibWAMyaP5VoCVzFCxRRDmAAiJ1x+WlixsWYHBpXxztClzJ9QOzGShLZo/K72HdhqGow4hStjLF2
OBREWSPPsqJjPxi92HjwAQx8hMOHCbkYdKs+T9H1EaPggkgk0i8iq7e5ppo/IcCnZ/TH4uzetwzY
w6GmyJ57SZLIrOX8ojTJwcBSHIwNQhzCDwtVzeQu2LWX93AS+L/dvvbW6Gx3zVRJ50rPoo8HA3QG
/xKeWNLc1LAynoY7Z2FP9tE4Sp6F3a7uWsXQ6vUKFXmgqUi1jZZn4Dgg5/znXmhDDYJCYLobdbut
d0KIAqwHnDlVbZct1+/7ES5nd/4TjRgkUwASesV1ZdrRV1CU6rk4TEi1BkZHIDXRp29GxOEaPosY
Vtcq4fVtjpt6bO7HKYHLHB8CpxkB/iCzyEYxAXf5TBSLOt7c8Ak507EswrzXFNmj/Z3Wyus5f1c1
fRN66NMGb8ODoj9MAnEiicyYabJsNlNYqZeV7o04bmHQObjRxmwnNqj1xyqCgeGYBNsUfdFQTV4r
a4HdS/6ZK16Ps2c7vJLoVCnNNElrn9uu7+G4PWD9kRjhPHRPEgvmkLeufPihw3Q2ZhJyk4cf20/8
d06/79Bv52EpVHB60S+kf1emM8Hhaf41Q7Qv9baJSn5QA+a5mp5wUtZiTuZeIhdULz5PVe0Fgl52
StNswZiZ8p4C0CDMu8565zWuG8jDe9Psbq53MoovXU/QmUk4Dp4LH8UJLyyjcJnZO/DS8RxEuT+O
YlgjnFZuZ76Q7Q2fXt0KgBizgvhwwaaoi76ZyFXkwikz2tHmLB9MfyilXEz60C+VKlXNBOASPgw0
aU7zjLOyqCk7qD5dD4awZGSSbjWQjNihnB6sW4keguiWxPgihR80/Hx8m787wsud3bups661piQz
EHb9n+uGhU2VnLdS7naLcy1fcvVW918t9rQL76p0qOzvyFI0ECQfgN24i2Te7ksBCkFsevBq6Yg9
aBtpRPUnEuIFuav9/GbF+dP7b7Y2JZ7w7IpQfYYurUbzoRdK+kv2XwzqSF4jq1TkcWYv+/pp7Dku
OZvuFWM3JdTzKVlnEb98PmBdE7XAqTpWB0P/Pz0794FlPDrfzRAbrDDm6AUsgr1ddy71MaX32zW0
CsuPLwsJW+ijrP0eiUL1+UX8SO/vOD8ROavEuUxlsnEg2uMwcONRpb9KVtbHmjQdSVpArFbtYPAz
l1Vy3XxoM86P2bU3iQEC7b95zgEYxSzYXoFp52nU+5FFwtD33RJm1EoZBFNGQLfr6fw5UrNsPLTi
5F5RGpzdhpd9TMgROdE1FtINZIDTr21V/W/qWdCPjvf1Kp2WepXLNl9xJNrWx/kycjBssOT5q1Fg
xp8m1gJpV/QFDawx134rZbRYdPJf/eDJyzKbgAOspxQzm/UFiNF1c1aJkCbqIMNj+zBXrZLWeQz4
yyrze1gdVKmjQuo+F6G5UR1wTbQksKOkvAypyq425cTUUvN+P9sa2QA0XjCvp40iEOTONA/ZiL3S
vSp5DPjR/obgGlgH6PPnk/UVI+PLdza4idb6ZPwB0n0F3jbow3fd6cXFLh56Lu18TQp5cIvhdfq/
Kvrp0aLKX1BiIr1SKDh+r3iyENvPhRMSKMcOQDFDof7ZnbnLqWSZuVTEmV42nBvkukRyIkk0x4Vc
8JAxQhpsRqBvRp7Hmcj5qdX3+hcVs19rzb+oPvTZytCcz4xd5NU9qyJabokJJOPJJzPuHNvhvPgW
WrS3gEzEly2SNd3IYy5EztWblgYREjHgoHdjesUdibKd+61DRpT9Qk6pTWflVOP1oDDpPEqWtt1R
y3jXmIn1IPOHzFao6W5pZEYv9OZZVP9v49FM3Z9e1vOSnM9HusPKD9NHAO+85DxafP2Cj52wvT69
6j0CGOmltp/+OBMz7bM+OP5cVhnUZW+MSz9gJyAnODflZCWNOLKT9KWDksesrkSf69p3pqPVDUZS
uFXSCChwEKJTKqRzKG7+QnKeyoLSW2K6R5mCSpmPqqT8JALs8DwEkRy1T0O2ya+giCkuQAUKQUl3
AUivLoeduRpCBSlDpPMT92NXSgCiLA/g/E+oX5dRHWk+/8BOakSnZUlQ9mwz3OYAVmvK+86Z1UJx
XJY5+E0rOqim5dQTjACRTx03+nJ0NIwtFy23bmHujex/4l1DmiZ1CRZKEFMmp5abjr6ocmKU3b0o
TJeI14QKLolR0cHwt2BobMVMY4GuwlT50RqyMHd46mB44vHokUyzkAiPgG+Yh6bS/86tA6s0jzFG
MbQWoq5xNRL8GngNdDt/sMxjI0tQtgWxWBEDUgF3R5J8alv9zlJgmwBr0Rlnt/ypy5Ax7UKxMq/4
4VeMBoh+k4q4wiXpGM7DF04BzVZD4GQ63kyHPXA3Ur66vzzq37Alw46FyNqEknUM10tpjaQamMn1
pIRe/psgtB87a02GZX3A6u7vM/wMXjRzkPcEfvu6mVC183i6G3Z6fcZMzZazUNttuMd6PBVYXkB/
hpt7nudGA4FAFr6oZ6vdt2xWYugKwEm43Y+MifTNSpzPlOS3DKAixq5BCnykznPP+wz22/7SRhaa
CgIp7H/iuFPOm0nCs3LMP6jAkgg4bZ+7t+WfrmkqHzNZeow+0XfJ+Dmhao+j+IUikl8btclapHEF
2VscLLRrh++kTpw0UDD3YLic2qDTD5HFsvToNqMeQRGMH942IJOJ17M4bJEO94MwHK45Q4eQ9hPd
QbN0Mb25NKBGvA+BYbH2btBXIA1skKeIplruk9+0qNzoD5dKlbqyr9zYCy+R2ia+ZJz9xC+Ykm4b
w/O2gU2fJGFMc5hyroMgZx7G3+bkjydFH1Z6TZlFpl0u8EZs1IxskVMkqCvaEnuuSaDf9T5jOOoK
wpPCnq5vvJ2d7+eq3010XqfFvNVHUs3lhAvV2bprL+Xg84lvELSZeyyenJgZLFXzuHpwAOai9zhR
FFaPTnLeg5cj/Ao/0bLXL1pm50pa4bBJHS8YVDl1nCGtLfC6R39lp+JMSpAFpST5gCNHHwRvjJje
uWedXbUgWCA4wZ10ABACrG/hVf8WWMPM87YAygc0YF//IcFWBScuI3WUl/h7wBxmNjhZMDnrGOzi
Wa+1bI0I13naMT0SuczjC6Sqw9uRSK8elJR+m7gWazupR5yKT4zrC2PGuNyGNJ4zjuXqbPp/iLlH
QHik7mRPPbMvJ95SqtBUruxHXmbq2l3vp/yz0AevojyZCqsbeWYIAWQaiBgLSiT7UHx6xCZe6iXI
+CEpG/fb9CRXvs89Q+vRUyMdp28uf6PakFa3e4+HLUGGeAR7KTFvGwXyE4ECMLZSsI2f/zDRoRdv
rYk3Sirphuv6UUTnFJ42etwOV5ZsGmCpGYm2vID22jugEpGRm5aZayKiRuLqGgkt4rN6GsRAhscf
JaQETg1XJe8vvUhgQ2lUrwCt6ymYMU9VioBauWawwvb4u/MP1RY5PutueBJN9OrDpyteBwCkSCpW
DFrfpU/XlwcZ16wLJx9qcV55jw6PXvyeYfip8VuBFhGWv+x7vH3E2vY5wWMokpRUWSgZJzVkNQIq
aYKX3WDNM5/2JcOqI3dunZECHY3WCmMTNHSf3G1j9+a1sOUvvqazGFmXl6KUi604/IBsEbmMhSwx
vD5uH2KYRFey2edIGhs1DNFl+DchJoKkMxmlGqEMoMu6fZxfJV2+Ht5DCUZs7WRq13VaZN4mF14M
Wc60lXIdbq1lTMCFzB30HoDYPfFvxXgJGfCQaftj5HANe3sJGXm/E20jmxwFvQpqggtfibFr43r6
i9muniO1Izs8uTwlAhymFhkugp3eNkfCDvefTe91no+VfON6g66S/xoEez/KUBjVNwNYatkwjwbu
K4EFRKcqIAdOC8QVUa5di0bJ3BsSCLZVDkETD0C57rYfBCeJdvdFYbqffB30qUZxZJKEW64vUqa7
vGtIAxUroAlmwlmUYRr24gSspW/utiNJon0ZaquEnneqYOn/P9US2DjCfGaPoOXEqOx2nogdnCzz
Z1qREgsGAkSkwcFPjtC5MzbkgnL3ICGIb6ZgE5Uqt5ihS0KtNSz2Z3pOv+pe/+m8puJ8rny9DofU
kXqSnCCHPBRF3CmVnbSN2xkF6+FRmntgL1YQIyuQRN/I1S+O9aHF4yDZBXLbwb3qOmLoxgcafUBt
tFtVxPm/0ij+GzemHyJ6BsDI9OXJXxM3rGNczpoKN4Nobr0HmJ/Ml34LO/gIi2/WHNGfHFEJdPoG
qYYBkl9UdoEieJ46cG3LmF2BNCi/um9pT2MPAozYLXc2i5ShGgXxSW0OL3vFJLcqOc9J+/nX6yxe
IrwHjiEe5al+2IANu2592UWjOdkQWY3BoDjWlq8IittpM+CeGgPqXw0iU3Oy1OjFo6bqgsryPog4
XtKFezZj46Yk9ishZTmpI6YL1Aj/LcUieGxopk/HSFbATq8cqU6LXQ+3DM+0R2Na4PAE1Xh7h5vF
My8TE4QtRo4eS1tUzzbZ5DjOhWBm2J+DTjxkp1uqi+j9azlsMSbfxvITP+QW4WNN3GG0RcRHgP/m
32DV1s9obvUzNTtar0dBvb/y9BtK7iAtc+Q/M33TpdyPB1WQHJpx33psbmlez9iLPJENxqmsVXY5
ZAY5hfRC/iXK/AiM5k0Fvn5bwLcCnHRnuFgh+FQ/ZtbIoQqhD9odBbkGB5A9Nr5upX5lTOyyIc7D
98PZff5LxanoMyYZ3ouBArASvrr9yUjIMmoPfibbjUZXFFohGwuUs30D1LRXFvyg9VbhO1Bz2wME
waAxsWfGAGyKjKGpEkIrYD4RRVjU8df1lPccUbwAcbHj2rAukecZq6GjMA/miNwSAM2liHXyjhKl
qb9LA6DnIUdDEt6uzvFNyLQEi6SJS4bMtXbUEVS72AVj9jbSSVpfqgr09vTfe4Dhmqghb3cLw1im
A3gUfafHuB9FAIkm1TW574GbvW0ZNN3c3fkorcGW1of4RS2lr1yc09NcJjZ9Oq8xXfx3gUHlKFBS
f1FZJ4RGk28Tbux3hPohSnGwJKdmRAukCUPnonCy+LUXUuHptUZ50osPRbu6RtfOBYyHb5iSYUPA
7dOg76ZyOTyCJvCjgXWmzqj3weDAU+pDnm3oGGmCgQ3DexRij0Nd/hnjnYXks8V4HHu7Z9Hl5D7Q
yc35Y9XjF3tpUyg8TcRPGhf6FuIr2/8TgQwkulzrhyVwKCXkCADziwrOWT6m45CP7lIzlDl17mVW
PW0OmnOUgecGdA4BmY846CW6qg8xewsXAolQbCyPJHvtb5/CGxPod0QXmuvNn8tN9qcOrZyz5rHn
qGzSguxAHzFaNmE3mGEmXS3P5oGHnWYczC/z0LjhzQOOtz8E+O27BvCIJGvU4uso/To4oVOzyXSR
R4rw2ceu8nA1FNQIL+x5oxgcyELJYf8g535Ntd+fckdckDJ8cey8hyKiq2oC+VvkLQcpPIMRc+S9
wCt77V5oweLV0E23xtC46js1gKpam6K2fDKkRi9ZdLy9QkinyxA5ZW28KajL3RtwinkwIq8QU48/
OqR6i0VNaCVXPoI02lQkK5BcbccFSlQ7MmPCA/ppROttdz315PKLVxF9SdMbp2ywEMbtyY5KAwHO
QhzvmSdOg7gWLJrNX9Rwe1JjWKq0N/rqrd+Jgu49xAKWAFXOdM+Q8/Y3MardejVpwYR7NMwhhzb9
A1ekK4xRnHVBblq/KEFBY/nItpeVyuNnx56AYKAoI0tbyy4S+/arTF4QEWH+24jXsJHi4kWvJDNE
5AgNpqH67KUjPhl+GXErqKOlu2JbyxQT57UaV4mfaQlCIzP+RGSOgXjx3wgGAAylsDwzySlCMHqR
MFdcKDCscaLKQ5oonb9EbuNHrObHUraEERe5+yMUkYlqLGzpdQhB3vlhsj4qP0IE2yY0EinSM/e3
tbvIi6Nt5gaEMgSHxJhecki5pb//yFlCz7sWioHiRKJNeY7kjiIXoHzqJP0Pa0su8IrJfSRQy08J
8wnbw9i2MDyUS5TmaSWVQak7M/EBuMDbWqJUcphScpCDJY3pw+hV8IuY/GfpK7b3XuKmyrPpdL0j
Xw6xTYLnQB+F9zcrF9QzMh1GiyhtBkkAXWzSMkVtFse6r0pxGR+OWCic6HnNuccZII19bIFNepvv
tbOgEIodQ7hp51ir7MjPhBUbavI9xFtSQrFJZxL/c7Pa0GR1Q6FLXg6qP0Juzs1nP5UJNf4l82nq
dHpzmSkLvq+ne87Fy3QZiYrJBmOScpEIXY4Tmefn2CLsJQt5H5DgbRR0xHxUlWo+RRmC+Q+/QtY1
2MWj5Fy+A2Wic8j5SH/lgYcUIoWN4Uq4VgeRFREBkcoEoebLi+CFFW+OsdchHVHQtJIbyuOcMGDY
mQ2l+cOK20y6Dlo5a8m/VDjBaYVh12umMbh3PHrnl8/dYR0MQz7XfApU3KNQHZPzVmaQBDalhFE+
cmqbV2Qqh3/7i9NZod60sEQWqQ+E0aUq0wri4yKP/jKTdAO295/FCw33Wu3ndCeBCQP/ZAbywF+L
zVlEI6yiTg1M70RE8w2xmeiT8Ur/6tcGk3YVXVQUaWC3q5WQDvVmZ/bSvT+N+8xSm1I9OmzoRLQv
aI8+0JEStR2iCB7fX0BGZfchFR5F3fuCM3r2QA+t91FVPqY7EOrXyDA22/f6MU4MI3IVN9E3VJBG
9YVDcLaRBdaUhzWPWLuI45b5z22nu+RxoiqAbALZQf+KVoEzZyeu14c0ztBkGtqlhadfHTHh0Igg
uwWXL3F/zqBovLSC47Ca24Oh43CgP9ocQX3VTM8bJ6X6WEuXaidbm1JndSMipdHw0mSTV/zO7kv7
VFOSZMAfn0bR/HtRG3AX1falTLXGzmxd8uQtF101tkPeI8RgODcBs/G+hI1NuWEojj0oVEgottRu
UyF5YKHmZoSuRDmh20WKt400/IEMqNhSkyEj1g8rTgWlDsn0b1gB1dqIHzvhOMtM28ZGDmS7FNhl
OgnD9nAoaV7Cd+MoNH/yajMBIegBUP9xYou5gD04wBVCeV1OIG/rDJwta7YdHBPCnM7T6dbIg1X/
GA6xA4tEYC1Ngg9GFxSnGXwL3JoVbQOirlPPPnUE6bG11ohlM0UkpSryfFhRf8VnixpzBUOwYnyf
yf/1qKqg3/p6o7QedpeMv2eEKvQFPXe1fFdErTVdkxGzMuhmawNlju+yGFgsUjaQmbt3SOvCFcpP
o8U9Jkp9r4xbyKu4ZwDcRkYDuP+mvPqiPYSVNB/TBGoQ5+bckt18RHmRoOonWOJJkWSDqA1eHdXe
DXrX5heu2VuhjdbzHQRJ/N63d5f+yv6hhUw+8z5EuqzaUHU9ojgBL8WZpWJYp8SwqGWdj/MGna0k
gXv+D2Mdcps54GbZr9iCCevx9gmlBDwBjtjjJAP2MWAp4fvI8+Zon4rs8ad8gBu/dUYHvqwn75I7
6UVnBlBw/8pC7a0ef0ZlclzMgAZAzpQ9HjRj3UP13q12ThE12OvURomX+ejF27Ku41G5yZyDfwDr
UrWdHBrKk3xarvTAv5wbTw4Nzl65az3/Jo8f+KkGNLNVzbxFi1XlyagAPoXC3KHSX9G6J89ty13G
o0MepS4fTHrlG084trkMqfc1lEF81Ewqv2QH+9A4dHUxcJvXQ31v7hxyxuxSD5rChcHSiO/iuQGp
PaRJoDSENaN27ri3y/PWkAhzjVnRs295YDS0tpxgyLfVe/wfO0irizlAVPgkXgY0Y7Eu9UydaXng
mhU2R04aRVNLnINsbRTQ1EpWSQycTLilP8qpnAmB3/Dxbi+gFEMyXtpZLBlO1/oqdwsNQoJ5OQaK
6m7p09jmHxhRcWC51MiIrKL60vuEnmer1qsr5/o469mtCaLdZRt6qULpT0hMK2M1LRu+XZhXpqy0
7ZHHl2aee5UnXeCIk7L4U/EJCS2ujwrTZunDzSDIObnYO6AO7BhpuKwEbaXc0Q8hynVAATOhAgtm
kScUSCXZ6TwkXQ5IeAktBm2KS2oygq7/5R63Uo0VmkQY5wsYmfYFtoRAuymzmpjsYgSpbjpepM6G
KieYB/2mnLpoHKmCIF9DGa5DTr1TagSTjNT1G7Cv7bBYbqGZxXYKsoos3mB2O9Mikp8q2LjDVHFt
pqBR4y8LNlZTXkXTPpRbgevMjGa0HtXFFtxnkCFiX2e9/FBtSgs3l0vuLkjI/n5yVJBMjA8vTckz
SaHxol4YQMt1+jJoL01xtNSKdfVc5XxHQ5ZKJ06epFBKW4pimPQ3VWcI6gFZpKo/XbIu8PpBIECr
xoZ0zls/DHevwe2zC/t7gKS9xiQlXlToEUYr/pr7lmB7/2nfeM3l3CMlysr1GydI43QNvz60n15d
HLe7vK/cs0JCZLzd4AAmDDaUVTAZNE4SR+BGiDApzBzKadtbIWRQRTrrraAAXV48SVhyTblm3Ieh
0bAbOpY+cdmSqhMwWX1xVWiamR47q7JhftCyWezcDZiSAka8kfsG6P5MQqDT3i5CTRSGl+DmSATP
EmDZ0RR0CrBWsZlvHGhZ1kb5UmopPO85qsoMMmvplVhxs7YFUpkaqAU1xbgoYFJHiEZT5UI0+bAJ
mG/077QYk/BbmmYHi2+3n1wD03UGBBSNXdi7UPxDs5EKlIHn7ZrMyjNnYCCfcpU8GhXgxTbaCpjA
oAEQBjctKQB33fdXpgwl4jWFvBntq2o6qeSQrhiFIJHaHmac2rIlt472yEtJHSanjkQ2uA1a1jD/
PJCCNvdQbhNaEdTiF7v6FaylA/0M/RC+XNFQU/bH98iJI7eGJZtnZOEI6yJSCbPoLkEWIuFx7sDa
Xjfvf7Qy5GZJTo2hOPNX9ZFb5YJWGWrmd8XGTllg5AUh/+FneskHZ5PlUhAIEWSEhjttjccoeKgX
OJpGGFxa2sN7anQbIrGRbDafjoJDiT/HDI8msuGKYTEzqiKAeXIZFxHRjGn60KnAvfjMxRiE91Fc
a4GWtTLRotNljLsnA68WNhSEzWP+BCP0fbVJD9cKzMIf6STlDrPbN8UiHmXW0TbLb9JmMhSUbH0X
JbYYV6lLEx3czTeS1hQZhdgtFIg5zhYf9kZZRArs/FVzXRTNi5K3L76hh6Hk0LLYQceVP0XAkrGC
1P0lUKEOS9Mvv9LFvn3+sH+hb/aoSZayrA5mW4u+GVfwAxRJ82lDvjGhxkwYf/0sgsehdBcG+X0d
fvwcUutLL8SBrvAQc1oLIRrqVSw0u+JYIExLd/XlP57lSwOQU9mvQ56QP5g2CXbW/o3C/jn13gtS
Zf69b8Lw5b+/tYyf1uaTQi3FMNyd9urS1iBO0ntVDTGPclVHrLOoJx34u9ViBpAaD4FtPwTnabjv
W0kdlkLjYbC0uC3+cBWbpLdLaVGWe76IvczkZxNz9jkYkoRTDQG9jwx0SwsFaE7F+AqY7QkNRrXP
rHJ0Lr/6G6DrXbaNXmQ68qJQjqffQY0jwKnYRxJXuLjjgSPoW83xtN4VworX/Je5AfYCCLV26JYJ
RRLJXc2IQgyn2Ab8B9Vs0DnQXh6dQ9mEZCsLX3A1A2mYwgH6LIK9qfdOqG5GBkYM3Ge4Luu126zA
10vR0auwzTmV8LRe8aaRTTplDHRr2Gex4h9xIOLIk2RXw2yMYaHYYNPH4wqq4hBeaFcdGAAenw3H
FYL+hMVbeZZJ0uaLDIeHCg2Z0M5kXNQsnaJZ+RQmBdZW4qFOD9Rh8HIsnU5Jjty79p9igqBEJtYL
ZwbIPidD9dRVQfTpRrhk1Z4uoW2D/3UUsinisgYqZPGLlN+baEiIoI7mLDsALnSjb/S2AKPhm82V
7cdBkLaiy4qgY/wrBrEJ2trtx/HbKi18s8lYbE7e/rs2ip+VOYPbOfhBfShhXc1V8OZhYCgFgp7a
yP0zhGH5it1D8/zMrB+YYKCizNkZ9RhknvYH+vgvg/pXpasgybhQx1j9MKeiWVhkh15LeJjj/l4F
WY0JruiH0A7Z64gfK3d/W/cMfeT3fGrtTPsNMVvnXkJA01g6peJp7Dkh71ngPvZn6v0tRIEwiu6k
/vhirXwaYCfgtnc02pn5l2fjKCBTFk5MqgOpN3FOeqsK+zJGPIOXLPxgvOQoNMGkQVVx9DWzrwP5
4RFZcG6eGuMNnuLro2nKiR3FqRnM9RFKxADurbxRJWDAsUmrBBTnMLdhJ1f0GEkgvoiw76b7MEr7
yHw5ewpFlzJikJ/UGRO5WXHqq9wz4eq+5+38BFIRx+SYHe/N4d9Prprai29oKKQlyPPglCD0nKoO
xJ6N76OH0M12JukY76W+kjT+dY4zYZJP8WTQT/Au8jYaCb5BRuchiduBpm42BPveYX0tikcgZq5z
pu6E0W1EZFh9aITk/wvDoboeQKP4upjXEv7tKGqpE8r2u4gC1wTti3kRfsVT5hT9IK2f/ZrcOqKV
oFR8WoW88E4U2oWjxx9jvFidrHjp3mGsvlk/3mmkEsXYpUGasraXyP3wu2Q09AbAeHrWInavk4eX
c3tq/VH6F3i5jF+kqpzkTOAVQkAbvFuxeI5gvaAiYELRrAnVniFW3RktEAaPdUAvsHiyHc3GOHyF
VoDM4Rj/0ZWuke+Dcb1E/aW+utoXTWYZHtfu6U/TBJSGNGLvgKYi8WcvRYZOi8webqAMnIzoM45A
Z0wBEkyPznP8jsBgDTdlMKv5AnpvpL/PU9DvHSEDnfB935sy/uggiz2G6/ejOppz6ZOjuiuRUlpX
JK7Vq2NDcjfQlfDTrbhZcrKLAYGWdP3wRr3+zBbBcoqdrCN8r7yNLKtkpprsd09bVQKU7el7mmUM
MTco4uEpDtsvV3p+RU1aEaXSCwlCZkCZ2E/hgMnsZsWY/5Vt0fcVdmI4Rf0acg1ox3yrdALEUK9U
sTKGiHQ4ubosBsNS3kBVd1FCLcGJS152YSf3hSkHdSKUEVpibRL16nq1Uw9YXrP7QJauVUpPH2cE
mj4Fbf4KZMzEnDXLSe1Wt2SFW3mYjFfcDufT/l4PB7fzZwhlPVfOFS2MIVydmmU8kSPKJ03TRI3/
Fjrrl3CliFYnGTjM1ZE4KWLGFlriniElKNP+H0a3hctuA5rAusoBmgf4yn8gUkr3agZfm2NOGrfF
XdxjeDsKKKoSumU32vjk9GUBw4KVWJ/Xd3gLgOYCDhmSDaqIMYLH50dXNzIOKv+7ORzETxf1DNXU
AGtALJPuscXvs8MX8EXz6lQ+VpgNwZa+YET9bdAiEK4LMc4WhNCZUsNOF06alpWuJUN2ByHUtGnd
D9mn//3W6RKyqzPBUmxWB4YfHFmsb7tH/65tcJQJCKuD/pOLBSbQ/50JQzHGaMQmYCqTWbQQtllT
1ImgaiQjgqRbEpyO8rME1gUoA698kWPJjMbgYmc0ucB7+A1HZ8gXbJTQGOWkgZ/jkiRJO4lz0XPg
GP7wtEPHzKkDRxddrAImLdrcXJqIpNxwB++MG6QQzX2nFYDnFJRouGYU1a8s0u4P0xDiK+xNUd0F
HfJncxSvDPQzjzKj+wzPR/H4ZdmVx1F81PQK6nbAAvHWr1VQ6bgOPCWY4JVxNQ9Y+mucxv+aoUFn
ZueGiLzYihZ2gLvri6LGbGfVFCMHTXV06dDP0qRcShlO85w+K7zUiUzx0q23vqcfXDBI1SSQuAQz
u+adUugCpJ1V/W96VWoPPrY+Yz2rjq2Bnb5Iq9hOOpB2vHOOE/FPqiyo3xdqqD6jnlgK3WHlDkaf
TH6EO5l0tnUnw3kjuyqgc+FyXg8O4ApeiyKTtR4pdRO9lrd/or8qwzYjkV5IsT/MTVXFxvQ6jNjc
Z6M1qAH8MqLEKdM8Sb80YqZMwKX01jV+yGY9vpiFwC08e8AS6NDFkzlBe2zV8Z2sS1RjgFbldHX0
M+7Q82UxrpHb8+NSEJLf4sCaQCtkp80U+MWRJiY35tdFvv8EwTqrKeqUNEMvVMWJMuIqtaHy2WTR
hI2zlOYd2rxOcRnIZBQqgueei57syXelEf6CsX0x5HCQ+qA6INh7M2w4U5u2UApHLJhEb/TUHy69
8eLXiCd3TZCFCZbdrbqS7jOVyYtSxBZCEHzip1ARJUpSWL0Mlxmb74R8rwF+NxxyXLLg0veOM27s
VeTdSAyvIJhGKDmmwS1MVICbL2QtH2uUxmfRSDf5Bj9xADsm7OPhzuQomBxpgm5uStwM00wGCXu7
3TArxhhDpJl0a/Nsjor7VLf9CZbg0JcrpaAAXe7bGONryrim0O7XinwFPstyhSZQxT6TnbWJ8whU
WLB9ZvoSIYPBzo02KwiMV+INdE14FEIO3sYJCmzJkL+U+M14Z2Ca4HEYE3mZKd9iNMYUHGf4mlAs
XXWP9/oVx1yhfj0qT4H0KANr19OYw8yUhs9YGqKcXWyV6440Att8mkYCoEQAp+KXU/pAQZltaRCu
0G5aGZWmYwYfBHFTOIhiurVV20acgffsoEamRvEcxWgd+PsDnBlfZlsZZIdL7GStIWzWA69sgooI
lKtVEj5p96bHOglSFvGLVy71B3KCEnPxz1s6sEHSAYI9bRtMPw472UY0QTIOYDxRhsm7MJ1s8im+
RtrHZu1H3De2xTSUnYmTpIdkxh94DCvSN2iWbpBesW2utHn1jOLqOEepaco75DaLpLSJN0TPOyo+
vlqiv9RfHJZG5oUtGTpLW7YeZmlW94gcXgU1rfLkA1pCeWYaxMpF2M1eFJYD6+MugHXemGz/Atl9
t5Q/uyUAKuH2g86W7He+veTd7HJLTEaUvNXWkag5IbloJazOD6vnswowUErru98gDLf5rsxJvD/E
44tNVaO2IUPxSWodL3CAqhTqHTsufWAUcG8ytVtnDg+ZuXnMWw8h5aBrfXmqVoRGQhz+6Mg5VfEp
+swLABXt829HiYbHI26OVpWk6R9C/1f+S9CI/M6U75DcDEVeOFQo0131Buc9RGIwUz84Nch2bIzy
4HcduZ4eWkJXlBxXw4hbdxSbnAYl1R9qmgEvam+xr01HS7AKzJTk6ZbIo4EyXEsvLsNy44AHeTLp
PgMj7GvBQLhFXtEpRRxqDtcwKAYQV+xOV5vI/ADQsvFr1DAlNejyBAB9X9fghGRFOlGhwEDp5LUv
8s89XeO2OjRCVRSLMxyRnYT2llxeGVVxa/ai4hav8fkG5UVmhWSp2noUB6l0JLF3lzdFOns++eZ0
nJ5PJPtnahkBJbm1PkZae665iCLUjHDz3xYtLWUSKFQ6lFY+n5Rwk3UKv9Uf6Hg8EeKDjRChYCDC
jVwFZsdV5LqAELCu+48B4tEpshsNYdtcO9lN+qFW39vIMTry5JvhpjGZurSRLXLxdFENceU0mr6y
PptrLC0BGZmjXBAsGkqMxr1BP3g5USbCsprx3zV35FxjI/d/UwfE53KhXUBRTx/Csr7F0Vj5W2gc
F4MV4k4KcHTL3cE+HOQ6V0f7Qvo/gyiRsLooliAiLfeRNtFEMAOWrSrHuH3HK9gANzooP6jT8J1B
ViZnOPi76xF8L2WqXg/ROFcxprhs3+uuFxcv5gQrxz1slapzF4PstnkSygoP+bnM2HORANElU0lE
KnhcWpQd+dHgjGZV4HxZ7+UnXbT2wgwYx3xTQBMBVhjSp0YUeaqgvL7Evb0aKZRcE2gMMijUOduF
o+VvlxCRtTyCZT5NBda0y3rzZyzi3l5/VU9mtF9KdW+Ty7JcQ2T0dbZk/llSzkhGXiFzvWyisEA4
75eHIJs8/ZYW5hSlaQFQbQAxHWIDk/xojlW40LDTKeDqa9ftKVwz7HlHH7ou3534QHlTVwIVmgV5
n8G3jZCM6To7GBcPGSTxLaV6J5ittT/1c40bQ6dj4WPLL9CpVecJSMAvFrGsfH3kywSYnRzg1Uhb
3ThnN5oQXfBzcHnHeLk1/ZUAa6R1Ko0qTIws2GNVcYh2ibgNK6m5/hRh9vNMMcgQfiSoQGOqJwKY
Z6vLw/JTADUH/5mWiiWX13qBz5DIj7JLsZQAhoiM0W/jVcwXTavCDBxUp7hPcg83RH7Dhk/GHy+C
O714Fy6rsQJbqvXYK7hGy/0JyR/uSwy3Z98jwJn5eJcr0H7zwqMRx01QhZdN6m7bEtrKRcAN9jAv
JJ5SCppSMLUMRxWYRL1zkMmwu8c+D3seFT5asykTz27O2ymDRMbDgeQPQRHacAOFyGjkQpLyxfZV
ZdXP0PBSk+Wx+rM26DMbIGW8VzqNcQDH+dViM+UOmy6sXlAa/fL11OMfxxWD+m/yypTvoqCz7PfD
Au5A4lLw3QC9c9lQNpP4e/W4aqq0RHDez/ZNc/ZZ7I3VYIWzEWR3xejXqHSZ6fGeJdy/EZCjvVTA
Ozd6EQQ2oy31jbq2ryz6QHKZGNMK7j3TTAqmZtP3RjmrkTB69lL9/43YxjNdqyT7qDuyGSbe6tMa
f5r3RouGsnkFOIIOgl70jGXeMOmL/VEJ7O9szWTbTxZ3xRtERcYzBKrhqX1E/s1jrfYV0T/3lyO0
TW7ImQo1meSiG64ImPaVhtghCcVKRDw/Co4IlYdTsxrRr3krfCZQg4WQMXtbQ/XPTKBoZGeh5903
asdia98ImnNcq2o9rh0Et9DmRY6D6lYWLHceponOyEhvMUk/xL/+oRUCx3MzjvkpAv9FBGAN0C8u
wDqk0ciX62e6iZLMANnItqc4AoAVIjEQJMS/3hDqqU9E8wsH+q1DkB56H2VpN0XRVrmTs6lN10BG
KmFXd0UYM1t7GtEDba36GQ16ZvcXGsEFwsbIfrhQ3Zl7Exyii2KRJLvL6s/j6OAo3FS1Hjpj6bP9
5zd07CPCLv14mLM0puRJ6xtqngLl+WDPpWvuIr5x1ZzOeSbXQQ2owmI8r+DHzFbJf7vy00o9aPZ5
dossv9Kczfr+b8J7i9kWosBjyFWzaKcTOuyxP1gyyJrygl/gs+isgLWp+5Cz6arxF6FZjN8QWzHq
KLkkL3m+qKNzIxPexA7dRxPXVYmP33pFTTMwvPz+9y9jB/1Retuz597zRzrYZobBlGWlJ75maRqZ
aheM38q/EFAQLz5WOl/93wwYZQi051NbWvzhzIgxfEvdgAAMkCTn0u6+4nLEYUNoHf5Hq714zLzl
tScYXLzcM6JjJxBpkq2DexIRRPk7pIDjnzD9vLkhhmh1W0SEknTgeX2M7vESzqbUbBHmB7Mdgxlv
MwkniagGd3N3Xj+pcJBINjOLvmsn5vt9xlAFIuPVtLYDHNYM3Yl4tiHNZK2jnDvtF9LsSvLRHg8M
JIFaFpWDWa7wplZK5NQa1lHt+cK7XtUn5Pz/3AoY/mz3gLotou6Torz3ItRyYIE0ryvjOgAKPA5v
8JHmuwHlqEIfHCp4i181LrtSOnfmqF+4VmearC3jLqMIF89/ySPQ5SMl4QPiVGk9pudZFmVq3xvS
4WbgmiP1xb0Tsev0vuyT3qoJLe9la2B5pTKKtwoAuvdwQYZF0DLBJnftgmboFLkRAjlWMfp69oV6
HhOguPNk6sbiV5Bxg9MOELqSMUrexwx4ujIETemkcc2+EWJYQ4EJLNqfTSSHAwguVeZPrmo40dHe
1lgXxqnLOh7zpklnibUmyTSr1+iqzUZf+pkru7ItjN0vf9Af6H3LBeU+UuYCHJXm3qefA+OpLUAP
jHSKGfbApPmRg2CmSV4VOA/j2tIrlt9b5mbZIRrGda+StE35ryQqH89BWcaebHTD8KqOYcJeM1rm
7SZULGQpr+DN3VolhKYeEFweA6saRXh8S5Uv5sK8XQCt5a0b3OiNsPgiSnKbSmbMPIxLX2rEHlcz
7OaDceC+GIDjUYTT24KShFKWya5E66SWrHsuiUcPTiqlrZ1mcox6oe2Zw9h4E1qgOI1+DwqM0e8v
6SbgBciu8niiX6v5QZpULWCQNO+2Hw9yrGXeTxYnG8GPKtTNGEQPdIq6PjFgzTGKj30Q0qJ3DfdW
XP3y8wkBDCAd/8GsYaFaZCVPgkCRTjiHWV0gpqeMktijCkgMPPfTybh5/Q0y1SYkW+MNMeGNSbJP
zNkEzx+c0JAvmZofin5pTfaCf25r0ORP70fEb7ivn4vohV3DJRABidYx40LrWMgTYZztIvtyXSpk
BKlxBWE3tg+gRqOIVbjr/Eprzsq18VWVJKPMH2ZXHwJ6axBILis1FbHx5LbrAFM6m22Sa1mNbose
f4aDEg5OxiY6FZ/uzYsqJllVvS1AxOOmtn7dB7ufcrNGyiLrlLuCRWx8V5zaMbRAvlLAsZ96IdSA
KM5Me+ys+DgwCoqijS5REkwYreadLNEO1fmD0mXd4U+h4AR+r+4NCySCsmaxdYt5az+HD8ONDK1n
Zs5G9NRJ1werVAyQYbCg4sfNy1WHezrloYhm5k5FaEENnC8XAFof62lGN+89CB0XaYkfmJm90SEA
d4r8vtMTvWW5bXG6nkAGPRwmyDT24Th4Xr2kQpc/zzY6VmbjhdbSFSu6TjtYGtkD3EOH+qXZYaBg
5mMkR/8fxp3vx0vtTa2YvC2kGu75ktUfGwzHsF4U5IuXQKpoudWriYrj5EWVoBXoXlRioxYja7rQ
oRey6Cr1v/W3onpO/jWPRHB43zNCg1+XL8CtJAQv5GYAgd+ZkzShGt36hp0lu/KeTdIYBGAy1m4j
4Aw5pXcW8zG19zYKxO5z3a1gbuDQUKUN78tjNyjaFoN3HZLeDNOIxOEfJn911E+ueT401WAQMGhy
W4n+VoBfg0QQ0Y8UUfUugOZlLWe1tGdWXFahWWSV2NT1PtUMZPxb1Un22XS6BKBrq41OFa+Uwm27
ol7LRNGl9XbFAuL+DvxhqI3/r7HDraKTLSNAcpHG0dtqGcGkWFQ3U2HKg0bGXt9ksg1rHfZ38VJq
nOXgixWc+IhXwtEQ/Lb+yEKA8/T4WxDT7/Pk/EJld6c8TakiJ14FsCnOSM5Cn8ptZbgfCOcsJLQw
i5RuXRDxhyOmLaLHHx7BU7Wob88FNAHuqMypqZ6dF6bi0sWF/kV5OAcTssI8NJASpXghobyb9Fw7
H/z1ytfeu5hnimP9RqjbFHwipJcpCTrdDSwRL+FqKrjojmTPTlDagP9hxX13UUlXzQv9h6AoOBsT
imP1MiumilIlQIAhi++5Rkps9bg4RBPk0jw8en3suFaGTFpeCQ0dmj8QUXrUzPdPrk0bk0iZbQ89
Mji+4RhfO33NGUue0M3WBJcueFKo/TA9wO4ynBxZv8G4l+sg9hPj5krc+p+fy/nwTF6HymkzZhP+
xBArgXMsKxLLi3RsY+FpaMPI1vd4aUlF8sIQ3t5fbzKeNaWUxb6hDlTlyejAOYVp2POR8CromPY3
ZbezRCwp6hlZ1w+spe88wjv8hT6yWGk+M3bcZQHWCx4274xOHzIt6BYxw3vjmupUPm0xMUQHaMkM
jSRekAJXTPWwiQ69BG/DhRyLVMHtJqGRvuwe5e3dcDFz4clKbCaymo992Api3Kj4qH8WT9Y7384k
8g74ZFIYJ7YYCseXE8aRuW20N2VoVLulz8llSHjMfbXVQy1HX1zKBmqWSxW5n0o3KV7pEkZrzhyc
AUvDi60558XCtHZyIneSDfGbTiuSoyh2RA/e+H+7hIon3w6inyc13xu8qkAXlqJbpw7JuuxoDu0H
/NJ2m9eH0macxKJVCu32qhCezm9s+XYDvGhxQ1eCWt3/nwr/FpeAObQHE4BxrnKZW4RHxllJJYSo
f9/q869rGJ4y+jaeTsufZPW9EQuXzUJR+dgPyR2udX+OiFTtX/oKXYRKn/pVexwHcIYRLV1dx4Gq
8ZHSFoQEjGuJ7nBMRLkJND+ohee014UDPIFySL9ThCKxr3/ITDJU15e6Rx8qUJ1QyfwDPNuJsx6g
HHLvaB+VbXC+NaF12M6tmWnudLN7APXep+hEmTaGeS3RiOv1MRE7n6Qft5D7c0GL3mgKlBnO1Mgp
Wma9Xdsx37jEiFw8/e+cUwbCZLjDFXLwsXHcZNkRz4Vq/Q0Y0nKDGHAXRza7lxhqHQ2PDE3SfNyb
+lFGKdHUp4g5uvfyCGddd88xeAdt3f92Sxo7YOH6e3wW6zOvY+oOWkVC58FwTL0rke4dn9N7nIdO
OgHt7uH1FUH4bixMB1MIsXE4ygEf3CbnjyB7gmhp0FvsVPn/wqvaXuHlzwpPY/wmv82CAxI9UKTA
9AOcyl91Uzz9tbVs3ObB8h8H2UZaqyTWJ5kNrSTm8xj2xWxrNLjxXgItG2Zm7NqtCORY6lGn51Sj
NyQ0Mth2SMwIDJspEGni/HAs/XlR7ZjUkFOFeLj+gXAuyVWeD3cdqHnCNmN6nmYiW4khPubNa00j
tGrOFNKPSHeFvb3lwqYNMNpwbwFcocmNUsQHBxYSDy8Z7Wai3DjVBTBdNY30pGlqr+3MevBeA+fO
deoIOb1drxVGh3b+HAF8UgsCR0gBrTA0i3Y0gFQ1Pur4gMpfFYUtn94sUl8eUlJAJRuYd8seBUXC
H08u+dGvyZug8ERtpwIasmF2UEAUkCq+R4uIDtmqXLab06bwIBxX0nzFdnMX9Sf/E9z8UZXnwZry
leZ49WY/+K7dmzLW8N8o2AHjYwVhSAa0Djan/v4CAiMZYwguoO7BlHmQ+ZfHzpLq/hYYxKrj1FGz
2jlolZnydKMicKh7H5rmTH3l4DZnIbBh6jfO3bgQDvq9Nb4PAii1zvIX/rhvc0KQ0e/uqvXe38Jn
qCeQBcnGFqSWhtjY/xhFMSVHIHuZ/RuGwwzgKALumzcjypKu44jVj6NG/PNvdNHaqFx3SqiBfVSN
mIOGDshNiXxxWzMR2iS8bKsYzPHQ2gZgx1PdCh1WeoOakbqYbV0Ce4bCFaR5M8LtwYdP2XBNsgK4
V/o90lfBNinQyTiud8OyZH+WM/us1Dt+qC3yfWGR/t/4I9zgwA6kfpZyuPbVA/ZChlytSIo3/Vjf
dqCGD3NOPnp3LDQNc8jthZaMW4eqLOgpspJbg12fuuV0eMKzGe7DuHCpE/r0OR7dv/40LFDAjld5
Koj19V1sHnzAZUt5Lbt4LrTyxU9LVmgDabOdHgIbotSBU7eH+nhksyF5SELIstDqLuTBi1KQdlbx
pSMKKKaT2EBDJNdFy/LCWi+Y/iLmgJTY4LkfqrlcmJEdW7pfCnJVnsOy30y4+tCTcmWLljEt/Qsl
xQF+sAt3dQm9bzHrLpiJale/tcjayT0tFVtPQl4X4Qq/f2yE8ESZodG8TzcwKhFnYCfzTURb60AN
TsOGXg+O9u0PKmvg46zDT3xEf/hYKqB8+w7PIEtxXiUDJCGeYeTExsdB5YptoSM67Qok+/RXRaFD
0RtRGdjUCBo3rk7A7Sd766FPgtEHKzgs8IFlAz+UQOPZC4D7R3lRxaHWGrPO7OiEYvEksXTndBUQ
WDCG8AjtDufJSYwDBzxM+vVmgd+BSIPHtbAggDdrQG2irIWMJYBGSlYlcTbo/wxcwkapl2q91InQ
CM7M0DKlMTGTYkjYx2tnq/T5peteZs8Gw1f84+GG+0yBbkG+DAxf6BM/zAe1Ct6gkfWt01bJdogQ
mzC8huCqZ2nayIsyXhvbHnHAbdFKfwcL4Y8VfZCA6eTc+f7td5h61GDidE7CrAWbDZM/SxaPlHIa
0qQqRID1+6NL+bNjxyopv44mVMagdy38HDsL/c+nt9COHVgCcDcBalyOG3BTkgfEIrA8oUv5/PCW
00B96hEy++bpWyLt/8tzMoRPWkohcia70VX8dABDg4pRVpYpcY5i/f7rtpJPUtOraxr9PkHOnbVK
117eP7L0y3971JUvdAvEekmZorep0gzpF2++LLQNA0xbm0rqfNQMSjma/2/KLewbqfqtp/FH8RmA
vIIZuiPb0RBolLtlUQzZilusmVNrWF9ofy9ug4H250xdG9jKR8hg/MJvjjhvUZpE+4ZbP892dsc8
pm60vqfG00Pm/K+HUwotDxhUmblRrTJJCMDRzs1u1V6l/D4eylAvgixAW7nwXinJpkHUsmTmb5X0
0kLT2uSE7leU2GNkZeEGqHNoZZ/0YN4BRQiL28szFPrdRXRt0Yej1cAYJ1lGruIaWyk+IllBApcw
UtZlSs3WcyAezONTq2DzmoM+V0NEGsXmfh5dHi5rPW+HrKGRvA2k3O33vpb6/vPdP/3SmlaXtqcZ
Nsv0XMCNbbWcCxo0MP5fGnGtop/FmgVS2H5QfM+cckPkj5909GkueqSZwcZBiIiOxDo2KlhIruhe
VJieJtpwibAwlnuPKJxsgJRNUxWhMVA2xcP9i6xVAfGvq5P1xpW9JHHuy07cDy9vIrLOKPUBBcxn
5vhcAiCmEv/UmIw0jYN7jGIDxUYsyWeI1BjQOP8XtsXGCYzXTUaeia7IKwVe4J44p/1ltIOpF3ly
bDoatujUcmBG+Ejzw5zGisRlyOjiMG1KU2BV9L3MtMcKrn767nrRR6rxGtVnq+DCZ/oCgT61YhUB
VcHa8pGbmYyNeoA0HJG5D07WgpRlA90AFKiaadYlqpCBPOaF2Iucl5PxMFkXDhR3/oRk3ZIWtRZR
1SBYYPeYRrhfzj/ZfhhbvvI6k5DMkTVLgNriFkmsptOuU5HZY5lO9cqf0f7RzGkyhyMi8JewVsiB
r3Bi3KWtQI939TQxz0DPhiUhNiPYIo1k2D62yyPmTe1N7RtLlYBLwpVVqQ/3up7n7SBurnhYRWxY
XaC2sJ2v+X+8tDtn5FnuacNnRG0kRX5kHPstNOjRELQB9SndK4Vk9xdBNQYHLt50/2/pKx2Wc0uM
O91Nn+hg2hyEEiPlyBr4QRX6kGRZv8LKK5r7guhHdl125O1t6iVvKnJFuA25kyiYcKxgKem6M8K6
oTIjVuJI106j5mHFq/90UDAkICQ4qROIcoskKH83xDNcgq6coX9t87UQb6nrd/pKQ6MTYXx65PFX
GEoxBuI3IBSAG7TVG70Tq+lo6D2QQ38t1Wtge97f5K1sKT+U1638joC6HMdZpjggNt5DL6CVqIO2
dh0Y444lUB4n/YDuUfA+0HVuyWxm+st+90d+I0aCw7SyFV/yJQRTS9/IH0iVtsYPhupRG/bdLN73
z3R9W7lG7ab4t/TJenQpTAarUd98AlC16lLhHd4ISZuIevvzSiLNG8NoK4lcKBRklK0nW2Fi73xT
ca7d+1KrztPyVy/0/IPnzkz3C1kOZQPjIaY0GeDJ1VT5vt2UDZ32lVHaxZxUhLlFmPvWCAXTV7Ef
AWMmBiE3AXed3Ta11ZVlrYh2edJE1mzYT+tSA5NYHtfDTPcpuaaBpX55neDqC6CmhMnFA7poV7PT
YSDlHviVkD2EWe5LCHl7IBSzHL5R6HCRqYxKIfZQZW9LvHVsrzWzClRe8LmZYFq6ZtXAxX/c9A71
58IIGdkSbYBivgh0lK7qQ0YBt3SBzAE4WlOL38dveN3PFoWpK+xFouV0ERa05S17gH45d6xMAxrZ
xC78BNTzqpiv1mRoHI36JRpXefzJFlu0yFBOSeXJBX63Lks7M6LeRX1KgfcVyz2JhVvgQaCVLMZj
b6I2ogVPGbiglVKPrK885En5evPove6VabwtAclRO5M4ljQ1uM1cdkiFOX1dpeUerS3M+v7NSQmO
gC915p/HJUW++vnzO/fpoIbgycovN65LSOP0lB/93iDUNRDkwIowQLeA+Z+I4J7VJItR008KCz5u
EtXplxBr8FxkJbFzY7DQ25h+bLgGuFEOv2p2Pw0juNA/me/3aga167YcR9xQ2TFaWydsgcJTSHCq
AuFoTygdyABeqvOBxC7ZnXTSAu1TSSv4jPOBLNTY7EsZ3s6K6PQyd9ARlXs1YZv1D08x6/644myN
2VYmMvNIduv6wgaiEKGCCKcVPBLCJwTsOBEUwoG6iYao/EC6HLWAkhWKTy559ZTmXT+k4pb/LfSh
yySf5vfhHqTBxBOANN6dg0mrsJF1p0FSgC7kQqjkBasJCLDs80awzdFupRMoXHFSpzG250fpbAcr
lheuwug2NEMOHzspqji8t3k+lgxruK0C6zlBLfWg6v4Jt0LD5I9GXo7HsNNksosXnzKvGThkefPk
aeRo9KaXB7CA++lxQnhWX0pqy1+S3JmZ4DWSa5e+AS0Io1IF8qaBiLIhG17+aprfHGoLDB85jN2S
lVRQb0zugydvj9aohsKzA4cJO3JbqbpfkaNjeJv05LsXT9ty5u/fmLsoYTvjWOzPBDpvhm32Kp0K
PrZaWwuwZqPh8LpHTaLk4ydJx9+pm6K+8wXlOeScKCJT1tEMIxAba2/BT3fU05xsO0pzXdgMUIdU
oh/mD9FZ3/9B7LYvlmFtK3sbtJP6dnMDlGdR2O+pGBXuCiVhgeQpW6MO10/YWlFmilmhIRlwu+l7
8s2yFJqkITFQLUOa/61tk7/HBEnC6s5+Xto9igXgkApqRVbSAlwUcVpCVGSW6AGkQwUBPFKSu9Sb
953w+QazJeqAX0I0gJOB+yrNRiaImmcq9V/HVy+nBh4H+zb1ntYxw7Hh7BPVmzdo+3b4qnMzZVQ7
BD4kcDqKMFCeOeCd/W4ItXqYh2QiAKtQe47sPPy1i+oNC8whGjnouWdaMYZuXmJ0EB3RBGHXP765
DMcunnKaoOPU1W/tXGJFuH5SOZEndfZ3oyuuTm6RR3TOVY2lIqZcXL08yUd0Q5HERCup6OyUsOty
g2FEKgSH+pYwWDZY39VMqQbdJLRbV6ELn1KkmIO48RgW9wo9Ov2A+17SHKTmBSlPbTsVxLn2/fEL
x3iJe5ipbTV8+yCQUAue1/VeE7lS2hiHGojuld4IDPuLOaHU5jdC0JZRhNZxgi24RA7mm51fTeXV
hms0FNO4zB7NhqsyQBjvEQ70u78ESJdJYXTh7wofixV3cTC69m4eVLxcKlgnXUbVnfUXa/Tn1esZ
RdMwLBSddpEvf7j96/RLQ5nFsn0DXiCVeTN9pcSWrYwXx+/bvdouhNNVWFWuG1vL093JQ+R5H8GH
u7ZhEM685jkWSKdoGsebtw0vbQlHs9XAQU4E9DMqwJclDp5R/F7lHdoMTh0mwHVK0I+n2BRN7zUE
o46ckC0VSJAC2ZBLhUC7obMqiNTtnPgRaVJNzDb0F3ckIHJoTzPhlr83rV8SOpQb2WeuFLEpJEa4
3sdwUXelMPW8ap4E38z2dziHsipyuyOE9qTe/Joz4lF6TQwnZiEQMeHg/pMGkLUk0k+NWsu+VkZI
b8FAceUjtH6cnW/Litz/oI+nEjMteDKI7sgdyIGu/BH7z3bikYDLgMXsUKM04LdZQy1mpkOBrLtk
muuiXIsOjWblkV3WiBuvI471luvt6O7yY+3l1stbVz9W/z/zodHAwX5d+UBmNfv0u9XdA55Fyvg3
r6rAZy5qzeHVw5PAHmdhUcA5tQECPFUwVkNzUSWeD7LMIIxDPKV3YhOSKbZUMrJb0W1pHKa1Jowk
mwFC4++D5QsRctZy1O3qtKb822UsMUqq0gwKTvZzLx35xSqIXVDmCnpTyGysdlyzPTRnULpRFh4t
rzcmrVNKKU4mQLIvJmJzVdayt0Rny7miU3EsorPk/rdo/hqct/jEhi4VwyEfDUbKsNqJl3UEXJgj
nEnBazRPmrX0c35TTNRgca+r3giKDPDJVJuE2eSCVjm44PKaVDbrteezydAR8kIPkRzXuCuiydp3
l3ONjxgsKyJnvTgrWiRL825Td7Wz5jG9J+htvpagkuCDaiw/o0dIyPUvKlM70BLW0dUp0rOd+UYP
1TAYECfWth5sFeeSGeJyKUo/B5Lp0bSIz8h77sNj9d4FkHrsvwQ9xP1Ba58JOiCSxpNpaP3Zr5d9
CXAhKEWt/uqnbmJ2llesO7ERfhcb0okvuPhZFgZ/lZvlIiH0hp+521ZsaDvOAgJeql9klvIURBrQ
XEMVbQx8Z4ZfiVeBMFf9kXx9gX3m/5yIM1ZLGCYnBtFGG4QUH3GETLIezwlgHd5Hz7O9FCX9X9a9
UL80PmeyFUGFbFEhOAW7TZI3ItN1/Z2fP/52f2+SyhHnA4VUVAhXyVRLLY+DN0tdWIQzjTIfaO8H
YGTan7B++zz5qoPAxx+Q1enpwfQMgA48zXW65AK5Sf60aX8gFNtlvJuiQbTq2JtSb+72KV3ZE97a
pjwEi2AdTIflrg7wOWI0cExuEsbHurOIsbgwdaucpwAI68tWY3SIJB8I1aMacZ0yoZY8bJSCorDK
5oXle/K1xezbv18YOQop5s3bjXjvT/VOPXxiMuTNtvMh+O/gLfsRzREbYiHQRByO6TPn1nzL2hF8
6ZtDNMlin+iqQBiDCr5MAIuf7Gf8e51KlkP1HFDD9ZIfT4yhdi27Egv5KT3vl1FC/fJyGSyFq/Zj
6QUJGOLsBgAeOS+kdGhaV/c8sl2E51TonfAqDK/PHi5E8ZWrcaygFvPZZ52H+vw5gR+N39eGsRUd
0/01S9HiQRtSFyjI39DGVq48TQo79VvjyB1H3AILLhmGvBwM/9Rrls9SzTvN8QtJI0Nh0Swj4IEe
QwR5Xi1IdbrO0f5F+4mrzDTckv/r0chPJpcRrKMhP26H1dlgOf0WiWezxbZRAohnUBALYzKqLB6g
wEyIhnP+NGqG5l7qmCZvdITGg6iVo2Q0jLSbxE+G9zaPKjuNBvaCZaWVe1BAZeNfY+eniHCkKN4H
o8DQK+pfmxpIv8C6iyYtZSVhsKwIyec/qtKG9dhPUMRuMrkceaigiPwhWirdicAiFdf0FtSM9xNA
ZwyGm1OtGtCWwAJjx1V2z9BuUtU2r3uAB6zgsqKDWonrTOo/JN92xfrrihMSBv1m+46kvW8mBKlB
P5ikKzeVhQdEbTNMDGsVyC/Y/xKlPPjm0tY6Vo6afrvmFBJKsMTb7hrPQFR0KJddncUA7a9JI01F
eIUzsqG2gi+gh87WSWDnO+MSM1+mZVGFtc1LgMNU5Ej+oY8TI/HgxyY7q7TL+8opobT6+kGfNY11
HlOLJcxnNhm6o1ExEVp+GMKWkuTIvWWwKXH9XRqW27cuni+gAeDx6UK9X00smNE/PRQ12WtATyIF
+m6pZ2Acd7wuQnfkR5GjXoRMdmt9GFZxJJniRpNPHKr53Ov+kdoyHVDwifi790cp+Fug/anZpv9t
edSphqnSpfMYmsIoHT0OStfFdGmpFH5EVQiz5haJ5WoDO0M5mykkeHOVbpLShXF5G7ZtQT25/JUd
iXgCy/WhgszGnXBGMIgRpSWU+g2wm1GgRK+SBhAtRdr7bwqNcpeNbLo1th9F+JfXL70j7MI8eZ9N
G0Pb99hxHlV/urTEncwcMYjyDwoein+Vr2EMg+OyRQYZ/0daaxd+GJQbCFhVQJBAIqxhwUuxx45f
KStS1yFTavam/0WSqtElbyW9YA227uldfwePOCUw/HNBLtUoieaUwSVtXUmGfJ3hIk58bZMYOw/b
eBheGn8X+lPJWFLXycjm4bLQKVBwFRqGHwsvUy2lsDRKGk34CgRZieXed1YJUY/va4LRKlI5A2ka
qyEtMCfor5BofeZif5YJUGl1Y6CftF3f5zW2g1/XEQazllV+2kwlKjSTwUUM79F6oQTZNCRy57Kw
ODKdEwEQhcGTgkcFR2EgnpTFKXDRRNdjHMbtnEfdhQgzcy+YkPI6y19IzjEKT0tzRRPnOcrkMIhJ
qxLdvDR+gfaRp2NLu7RcTlOQotOQe+F+6bokyzjXm0877wSx9l1pWCQFzXnC1kZGgXTJ/Lx8Znq6
DPVLr4MaUJyYABPWDogTYSJgPcwalJN+gx2PY7eFUzc610U9oCJfjXh+AtzlEJv6+OAzeyy1IUS/
P1OncP46W4sfuPz2r7j6RTpp41963TuVXUIN/5EgRWULnVbUr9JwbAmWlET2CI2eWPnO5UGyO99H
5KagSz98oKICO1Mo7izT4FnrSR2WXmuq1yApMwKcj2F8kQ72x2EHcAQ+ak2B5qgFjH+9/tz82LPL
vsxwpJHgMsUklNWXtWRCgr4MuLfgfnnE1m7/2u7gQ+gwlk2xy7KpCWRe12qPZDOLlvLAcAOgZ76J
J4hjSxFRSOGdGQga2HLd6fQBi8qmTOAAgh3DmNUTYuriFkb1/U1yuCHXK/rJVsQ2j7IvG0w6EnQI
2YwbJROkIwCxA+IUye98NNcBvDI1GPTCzmFA2HQon6GidFq3mcMalPcD87VBUgrDVZHy0B4EuHdv
CFLxVK+6yBDHV5aciX/DIe5H9Nu/lSFtZDFBS8ntLgDXgLc0Z34Vb/o+3mx/TTCDgYt9VQM3abMP
l7Er7wbPTAeHcpGuiHXzJapBXN4hk0ysxfP/dRPmQlje1BFZ2JMZhsqPEKbiMryLsGmJAgTwfQpT
xK+NGKaANcPpX/455IPAY2moP/2diQ2TQ+p6ll11JPCnFNa6sY/v9xhzh41tlMd+wNzOMUuNO3cS
gj6mxHe5pTHmT8/BXIM1KQFXJM0Z7Q02GXWSWMbolsDEgPB4ZgdoCVpYerLPA1kDN4u22HSZnT16
eb7lo19ISyQxBifD2FfOaboNB/1k+4hRS3IoK2napCPo4ZJur9VaqdPrngpW9hajzGL+DktRnC8g
WJomg/5BOR49jiuq8Mpz5s/RT59h361T6Qk4eSy72Hdn1BvfbffHPMr56MoSZBqEekwUFPV5ehlF
UC9Y3EsIjHKwqTMlsUX+DMu/7D2zleiEUerhTdutb9SVXcM9CGywHwEy7ZQC/cA/+G/TUH+4Kr+T
h3HQp9f/V8zgJXwZS+zmvftZ6h2lkSgjvHL18oxxOk34/iaB2MHOZwxmUFJkidj4YVa9SVhEN5bl
ymB41kdkMYbk7jS/Its+jTELnK+cLen8IJ1kHjLeLhCf8RD1ALNv17do+W1vE1T3CRnxfv/j2bZo
2Op0I1yALu71Bk+ox2b0xjRmuz4ABP5zx9PkqFuFGmmHCzboE3Q07SzzZ+gRwmpeMjun1TgdaC+N
nuFBveQRdvkEq1JQe4OWRMVuVU4G0zTqUDgiXXc0Ub0HcC+ytw7rJDC/k0XhlTcj522tbHeWjfa8
xbkJ0ELf0WZKUPhFQxcnd1GAfaQ9LWlthRCTEYNjL5VmondfwMniJl6C3ydp4xyY0lG+zr7eUjsi
Z0PB0yOyEZu9PGWBwA3zzMNf4SV3GAovdovQnoCx5IItz6vOsfFbTtjvILCLIP4c/Z+T59i9zzUP
26Lfh8QiBvFFJk30IE9NgOUZoP2bPtfnfLh6tIzcjJFX1ilzB5pssdJMWio4b42stnETKWFwH82L
T3oZ6GuYWH7KrRbiHz5RkLo3d2GDBvADVKjZUW6jGUpgTtEa/bujkR64hPUmsb1YA5VM4uUpkeOv
SwSjSEmsO4siyTqzs4lvfTAvbxqBylOjtYiL/om1CEPbEOn2Rcig9yAiyET408GKDfGDrxOprHRs
06tn62uWP9T0xfrp4L9HOmEn91pRlXj9tIxkYo1NIfm/g/DiAX4utuqC2ii4fNr0QTqr0Zjgb9G+
t7pso6nfwcOkNMSzijghvnUOWNbjZJgXZP7pKJUxPdD+f28VUB876APoX9O9F5rt3hIOcHwSW0lU
92xh2nW0G3hVWLZbod1syXLJ7GhDXryS6kqBMgH5RLHjWB3u5WvbbQqP8nUMIVqsUiIVOHlFR9rj
j7D9S6PGEbyFOVo6GWe6CxNAa3ConNv7Z/R6dXlm6i7uWEwd6X0eUZ9Lw/Xlir89qbvUJ+iT6ZJ1
Nv2yWg7qFLq+G1j87WjzSGNNBh6H14o3WHDvWH4wtKsxa9ex56AwugbFsGanv+iQoJXcgrLlrto5
35xYZ7v7LTeB6YrII5YIF1HKdfO0JRxMTMLwC8QH5QH1UfhxtDj/oEsk0QUeWRvhBBjFEcw3KGu7
/CeHx4Nppf3E9vA1p8IGpW5bZnBux3HCLSHXhef4UUla3PKLmUxyoB/COj+9F3+0kHt/uHq6vPze
ZiZOkhDOWv+IFrhn7uFeA8HMzYu4Hi4c0MvRDQfOoydR8537cmwOQVBvz/5iifth1UfhAjzLk5XT
KU7CByIi1y1Go+MevzY5PPhRmMBgchamLtrlCNmTd44yblFC57sqCMWw80Y3nsDUHMC/8zTALLoK
y2k5yG8NcJwbu0VoQsXU0J20/TBoTCMHuYVjN1m3Y7XOsfSkJS8DsQQSz0AYQznOMbv3hy6T/h4n
nlRdEAwb53znXI4XpVky6vU2clZuNsE25MFyywzvHh26jfQwTLAeZsA+zaETUY/Wk5KsaSSJkmDc
HuiAemxU3YbtlvUcfaLIGAJHqjaolL7JC0YSjPzNX99H+72i8bmh7Zthtoxm/ddYldtJlgWun2GE
cATiTfRxPt8Qcag7uWp/Qdq1Kql9mm2vMRvRcPkWqXWqWUqpj18WgpkeXGhJAmouyyoFcjsZN1mm
dqw1B6hiWLnbfBBjMbRE6yiscSCqrtRKBCPMhfSb3X+9MAdjXUUcHiZ3k9eKAOaifjSxSB2A+c8y
xH13dfiz7beJPp06UY/6cZjC0GOicScDaTTg+f9DDfQXobTNdbf616efW7Ig8zhCF1v1evQLZnOX
TCKJUpZKxqmSVB1xAI/UKn4BrS5QwSVUsvvHLLEhOoifLnjSAqiuEzahPCM7FlzMgSNK0Bq8ZWsR
xCNrwjWvm9SJQ91l4hwTgtLlptxKhf3h/7Rkk0XHL35fwmMpo1JFIt2IpkiijfLp6q8ml4Jxua+M
mv8QfpouzY/J6WQtpFR1UbbkdT6u06FBziGQ9QCgubhlTUynbPkCJ0unKWWlArbc1luUEdstc+s2
CWVmZMhg1VNrrtYmE8xDz2R72BlPwpRG4WqKat0xva5qxck2wEBChaoa8HAGZivymhQ9WTmpgg0r
ebFPbK87g/KzgdroN23LLMiiz1zCFpZVGFvnNo2hBAchugA+jsm1HSOFQAFZZCiK9uKf1WZ7O6/R
GJYjupHa/gWXF5Tb8W5ttwqNyrWWUf52ULi6GJzlX04/Jos3KVWvO4iLJmR0aAQZ5jyf4uuBIvM7
0Gq5N3GsnxxUjoxMAcKOnxef2E1hc0ozDTZj7GMP6KtUooM22ZK0gqhrNHFMpjpvNkSlmLckKcaa
pIMP/eYfPBcSxl127vGihhf06vDLGFUC/EuoymGQSx5tq8pVYvvgDqISb0+tlbBdHPBh6ifvOsSO
hHrz5g+X3FXcTZh8YX/2H6Anq/utlG1+QbViXnbgGWXEz7T6ej/LXvFgzmnqy9unZ/jPLZpHZnpm
vcdPNcembwRUA9mMc/00/SbnBr8Zkk+Ba2lt1K5hbQ4dZ17JMlkAIA6rUqAB5py7IjGZ2lHTMK20
EptOdSQXxaE8GTMx+6QGRXCQVnnLmiO4CwFxO/dPSRo3C9nPjPJ6g3j16ijg3cxb4/cTgzoRTZcy
Le1XCRypY/hM+A44UmsD1q03/X6TmBGQhjqEShExCRsDl59XJRe38e4i83pFdfUVeMkSCgNUTcav
/dMDQ+cM+7YmbRENOm7QnP7ZgrQZCUrBzpARXttU8U0wQIItkv031VqPD0vt2cvLFDTTIdiD5iXu
MWIngx6NTv/+RDeS3Um44dLoBlpJb8Xcsi7YfWt0OSp/BYpiZKPWXeU7sWfFWK/BIApunUXY/x6Z
1Y+0YbylCEGN4/Ft5xcau2Ff8NFb2ke/TY60blSjTI20NZkDTcczsZd6axamtdiPuNuzSblWaeAN
p3zll3QPs/T1n7wrWkv6dUZkyT6eht5mlpJKYVUp1lfHRawxSG7Ank8hpreF5yrgvDal8T+3tIPS
To3CI9PtEfMybJB+6xJrfd40HX58bCHHtBxrVvtzBnpkgQofUdbqD0ptgwcnm6N9eWILEg+LzDIN
Df0MPBAmZsOocCfyz69rtZ7WbYm6sGJDhcnqoWQhOGj6j/uIDuNGpW1J8nNK7oJ5KVlC9CYER37i
hDzow/3o9PDUZlWMpK/9sF5hfMFNoaCHU9lTN0NyNZX47eOam+MJ4otPf1FfE3tSqRtfYKbu0LFx
QRjpRIyDDU2enBr3bpf1VFH+pHfF3BNcMKc2xiTV2GYHcNwJhgzd5/cA6xr5s7zW1BW/fTchmUBP
YkQBURuKlKLY4bzk1/BLnQvLWnBW0tlK4QmB/42ySfpNJ9ITei93hLKsQvt8iRAjIyse893QLByw
jcvlv8xkkmi5tu+1T9pR1/N3K2qr/FW3hFFZO+5vMA71QyV6xpt8kv35lXAadl7NvUXwmauCKtJD
2131Zh7eqMsbznHb/ktME3y6CY6ljYSVL5OOC205w1MpJmX214DLupyIHgCOBOIVpUmO/ofulEjb
vrTYvk9mMsMfiLAO8JHIafR2vZivEFv/vjOxB0sD+o7HDZ7kHb1XSV3lOEuThgrgakqF5XC/qwwx
a3qv362Vuo7DhOQ+KR/T72EsC6MDNgLdlcObKGU2zsH/TURUR8dBD+w5NJr/EaFNWWMUZ0K/Irbo
3GNgI7X0nf/ognHovc+NYWGYh0wSshdQkHmv64Xhvv7sSKu7GQitWXZwrf/1KFINStCq6vM58rqS
e5AloGzm7DFxwVWpuSyMMYw4tLet/T8hPEr0byAIOmqQLu00Ub/3dt/Q7hWsPjRtM2w16gxEtRHj
wRafqxPawKvWEAQHNL0L5Hfj08YIyvfoKnW5NbjLogBuUeMXiSU83KE60mb7ItA3t4OPb29uQKaj
eXFSa8ZsWNMQ5/kRSwvkJ6uR9S6aYLusT19DkFkoXNsj1BOZ6FDGhj0hQ8YfGvaCLWhMRZ6IQwAE
gNoTGbQvvPYvYkpJP7WO/rCejJh/v5025vPav820ELo6M1TaasNSoidmaMeq1o4Ec3+8hzIiJNqe
YoEHS5aeRyxdNEiEtWySUc3ImJYgd8FLQRIGPjk32o6sR2yrfl0968I5vO+iYWHRVs3ci6pLnLJ8
cA4qZM16T03P4NyahOsxRP+6gEMDcb3bF6KSrKEz78Pt+uibMEDE84EpfF9gSY0Ydzl6dKnxq/Oa
C85YJpq5VXtq8mGtgwEQMlTul9L2V3HFbw8ca4WBglmfr17/bkwZbckf6wQU8R20nCfqcnk78mO7
yCLek6CxVRUZoE/jPrD8QcrVloxSt8kfW2MppksnuBGos+Elk4jkMZGN05aHjdFaE7wcJ1bqmwrp
vE74htSjkk2PinGX+4CkykXqMLCAFeAibOBrmG6+hhQbI2TmZdG9UmFKbpx2Fkt0r1JzB5C8G6QV
k0CmnvJ/EF08N/+hyo1GcoUQysyeY2vlHZ5NGHbi5nGh+cdiXljEsRyxsw+vSUJPs+XvYeeWgtZr
TdY1gf9oEzUe8IqeQsUNv5THx/qHhydopLZ38xpasV/gdzoNlO2tg87xhoCfyaNupuVGdhRrzOfd
7UwsxfWmuyHlL5UufW8fVBPYNY5+W4zQt1flSsaOUkIpOHRdZg+bPGFrEkJ+gcfSPQiOy1U6Szb5
v2oV/K9bzQ1QR7/nv1KHlKNpXQWVYBzIKmD77pl5diDVb+ObFpQL0lu0n5yJeXbXEBzBXvlHabVE
22FpQSLbSVaq+NdGixSgcx9CJHeS/aATcLlv+oM8fWnPXhP26DmTLZoUvtWY+7xCtlq8m8ALEn3P
jgsWfaM7D11ZxhR+E9r7T7H1HIXEVwZ7CZqzPDqVG1sL015++7Az248d1JieJXGBJ3890tos+en5
Ji2hFEhE0z/wMyzEzvCBLSeUBRWe8p4uCL98s4xDwsF0KXaqsEXeZov6Ex8DH+ajmJ1SuyCCkF8n
+zWofLq2WY6xqT/RXa//mgdkRDT2MjvMReIF7kdvugDVUk035mHPWermT2R6HTaXc5h3mNCu1aR4
GMiCVraY0o3KbvyBemurzaQRvaPMPpQvO1cp5/X1K1eIQEFbnYkEmQzn7j/OfeYX4d4259qnV/7Q
FcHfY9qVjmzmUAR2+4VzK2S5VW4Gc8BhmE8R25LuRiFjQdVj1yQs1j90LKV3Gg9ZDsPKfrFUmX/H
6Ty9gyk7TFfN7fmcJZDwZAGHmQWbdooAr8E2Pjh8hX1JhSBNbhnrp3qpQhTj7oo8myBcZenW3Pca
7Xg+k58MZ1UG6411/9zwd36j1ft2lhKfXFvETM47EZH1qlWxYlprgEMyj3d9mru0b+gK0ebN4zRa
lrJL9zsv1KWoY5G9v2V0nZJd3DfNQMB8/CETijkyzSsIMBM6evi4V5SoHuPHVbOsgbYaandnI0bg
S7AShBkdbImWi/uvVd+qEmodsFV4z32LSokXudnUY9rDRajgzII1iHz3j5d3VUAVkLuZsxJsGu2/
pi8evGYrfTW4Ob5eu8uLVqRsNSw4ptKGgHoBydUgF7pMUr6kamq5AjgbSEnE764YZME5bUHV1/6v
TRSUuTNhfefweUN2qPm8O1V9qaQZvHY6qx14svCdFeqXbN+OF31npjtDD1kgigwExQIhSPrbLiUO
q8tBN3TdT1Fl4EQYZ3jYAbS1/xnuWtlw9R+Avmqwj6C9m/pDpt+ALHY3jSS1vKczmSXVOOHO61mo
AyrAXh4W6SpNqw2pQ9g6qsaTt77DgkaPTAndnrI4jiPKk5oI4QSXtDjlIcipUsrCsM0nLxY/GTVz
CNC3iOk8yV7dePwu1FxyO7/Tdr89SSxzz/L5aOqjSxTKOp9CFK5h626DtgAamw8yXhiiRs11Byxk
bW1iGZhFMng+RtQ/4LdXCThwKgWIXimbSydeCB3KiGaJNGzSUXMO5gB6ivQ+k3F3kZy6NJZokQ+a
z4OnWI7gHVvkz2z1R7WIKxLklF2nalwoRUdKn0BoCBFz7+IaLV8qjAH53fbF7zXLARqHm14akVvd
DI+QF7gHrGpeqH0ICXahZTgBmeBVsP/DoEEnBNMORuljWHMjVETzhNTps2zy2mzpP7i6HdNpEh0q
aEA2mijQetjPtKyk1tzQTkR5jULNePxzkSP6CesABhxBGVo3vGvP+LGpp/5/rKXP0yLpJAdqhSg5
bMFZBJF7DlOrWM4cdU5RzouL/X4OgbdGCcqPVqb7/adATwbzyzmjQlKGtnylXKspndu0jJa8demS
1Mh9ORaZTnEKR075D5i6LbDvhpyzxwhfbqW80icXdqG01qIjoQoVLFm4AoEO9XZHq2oZrDVqFypp
PipLNAY2XPkwRx43a2FEFtVg5KsJTCNRFAUbxNFkw1wfrzoyP+flj/OVMei/ohsz7pa99uZc2yUm
cQhsjgmiIMQhAIyh555WZor1qYBuptCmkNlqyrDibpFSlVu/ln9WO9cJKrj+6zL/g3cWIYsRZd4H
rHbhfOy4BzUsvd33JDlGU/oYFPeGhzTuWfYklMWSyz+H/tcRdPDlzpMX7JX/NmAz4iwKyu1cYcq4
xMeb9JKGWHTcRusGT3wzPwJuvqsj76cIzRrrTvsAkccdKvlL3l4OFBBTifpPcr34xWYIJlLfZLhM
hky0pd3k3blAzRbaOtgN9ixXaJ+PVEmI+yk8zm/CQq/eSO7kZBINEGxceqVRg5ApCs5Zx8UJTW7M
iN2KDP1ILVYk80hZyVyvRs5OPp8+KzUv824y0B42lU/NBMC7kn1zJXHdpvceomVw4ckPlEiFsSFA
Gi1xGhKVjbx9hDlozNHlPSlUj4+25RhXJNiCApohP+M/xVSYnvqLBsP1mZzLBkKXd69LbitXq9q+
DJUgEiCUdXZ5MTKezrlO3cIULkulM++9e77PxyJNI98WuN66iQ7p+k0lMbVcIbrZN/FCIBg1CVEq
ykV+vid2Y3Z395dRl0b0tWJNQvMmaoI1XfWbSOk1o3N0CDt/s+/gZmUYYVuh1EkmNSUmFMCi+5ON
flhMrmQ3VHgSc+o0W0F+dMPCzdrzfN3hDY1rlvINGnoZtdJ30mvXVPdSFeGnVL7Gk8OuxGTJq9ox
jMSv3La4gmWBOpzgV8AuCA8To6NZIoLV5tnraQeKI+qb02PgrGl6AVMP4xA+rjU6a/e4wkI740E/
KzAeluLJfSxzMkAaWulW1kd6RDI7OUGVCO/i+k2npl8gZ5lSeV3wDQhHJQvSRZ1RK1Q7izcm7RBH
TrRGlODVULo/cO0PxZ5rLGJBEBCqte2ZPcQjXuUflTjEQTUjlvw9PoR/9cLHhHf0tMoh6Qhniedr
C53XulcWgq/DstztKtJxuEh3j6d1djxNIFe68Rjjs8NNbURmqrNupT9RK1QHAA3zyLne+NRB23n6
/On8FsuZhsiZ9Qw7K45TqycDMkHblsXhbZOj/LpbCBdJ5h02VSW5AJHthKdWiDnB8tHElwdNjYNb
cphHndQoN0iwyFgs6edsDYNsHv45jt/97JPtXgF/2MRjN1EOoU1nsNtXykKX9OPghKL1e+vLIy97
nY/YWNkfmZGPVqXzW6Y8FoiAl4bkjWiN2qvkEf0tl97EqbGFgRvT8y2pTDh8inzf+jEglMuXF/74
1jpixJ3v029A1gwyli+hg2YrYuyxl+gLyOSNMiIrzzGMj10fiqUINo9SM5er3bSdVEiUgWGnnnTk
TxXk2OiqR2lk+OlUMBE9haBCl4Q63zYOBQeTW5XHgjS81kyLxtRBRaSCBg3NdSamXuKMZuDDNWxH
WHa/xNEvkxD5SjSnRi6K5n3wpSa492+WKz2sIOd06gYpxfquUq6Jv8BYeEVnZfw03fgPPcyxLbH1
9yASsHovhf441yLVn8W4ZRxevcfTRiaTgj4HTQs5SoRD6gjAwxv7LfB58cT3tuBi9DmBdmdfwlov
2QynQCF3SxqywztndsuqvVnTdIpByalje5FVAIJWCl61chBN/fUpY5i8VYfhBPeouM1lQ2ff5I5n
kjZmHanHM+fmY/XVH6KaIQNqw6n2Rlx06PRTvR/bWVsc1GSqTreU7K+Oq45UZ7S3ffMcerowhP4o
MsFE/85uBZjdo8VEVqO+X2VYiqd1dVTuLKzo9NiB9VFu0em+ANTknH4SQUw/s4DWXUL6FR1mjhcJ
YiJ2EsX/3vd9C15ko+sFsuyWmQiAS+14Gy1oARPvNxLTbzEIM8RJ0GTYP5k/kt4PTHsGcu9u6iMD
Nuk89pvvu1nshPl+dSZmC7wK677TrA6zLRmNqPvX4FhEDUSH6sQTHItb342/4LmuxSMgefX1jwYD
faHmlJK07cuKMc42l90Pl0kg1VaLI0DeK+R8IV7OYWjAaLBtejhdC3rSgPagcDG4GOykQz/KSPux
8hnqYSEJSMxPhyObA0DtH4ONhhJKmtBoaPSSq40TvE83I8yfpkBo/+iauHsPLxRhCUWcMM0MblkH
bOspl8UOmBNCObmvatyWMYyqTCWnsdhHCG70yXPZy2dvmPCYnxSmyE9JfMtdWbyrlxqqPwZnbYbJ
6fzbKxjzhBNtS+Yufmuvl2f9cAa3UVzOxk6LFR4EtWmsAdsvDEGr5AjOC6fTSXb60cmEwYmb9PHx
27CVnlKuI0Ub17YGiBeRT0mDFJg8qy6fQ2n7XHIFJy+hIoc6Shn1hIu/GlrDv3SOcNFe1cOsDQES
IVI4CW2VqOUSV0FJb+/VAfnMW5lovyQcFF07tHf53iJOFYsboU0PqFvHF/2j4FgkT3WoJneg6Chm
6ieaTvcJs7ox+rsfEJ89EFSF/V4GgtkEb4e1qPQ5RCVT26wyXcQsg1+D8W9h2Z4qUTpoypHFx/ji
1mDxcfXuc/D6kQWdfKySHLjHyvQ3k1rZmHvEV4IelTSKCmPethSM+gB/xBMA1pTdYECbXyxkAorG
uSCmDFvOrLMrT3WEI2WVrKWtP/9qgDTfnvQu+jWOivt7BHdTiay19XlGzdIVy894qhVdTeVxOI9x
AWWd7ku9PwEslNjfiUBBF0Yupcz19exTxyjtGpuzL73ifqJEuOG8WtUmV3pnou5Z+adWijuQzV5Z
7X+h3s52TtDZprvUpeaGxv5/Vl9ZhBaZiCOIj56s3EAhJY+ImWN+lRNoTxcu8PK4hrV9U3Tv+ysd
gYiCL4T2sasuP4oqvNYl8nXkpOjej7aop384iTVXuMxI/8aEREX0F+cnb1CwQxc9ULOovgjOXMmC
WmPEfRf2KCse6DKtXy4qRcwAkwvNkqU5De/GdbD91HzIG7bC/TFUuJd8jcgk4HJt9h59JAuRoSGF
WIGJjXnJmXtSjyYjVUyoPbdQ2PBVZCclqHoga2FUPTNksEju5ExwDS4qRmJFSHc6LrhGKm+j2zYJ
qwHxLL/mVxyKEQt9hRoqT9XvOxbJFOKPTmNMnynKiGjg2f7w1irL+OnffcHP4AYq33G3w9d7T6xz
E7j9yfqUn/H6gsREZaYt9w6+fKRLBRJeNZ+ZtQg7odRsCHX5OlJxr2+7Okfk5F5QtDqvamlSRT66
8w5JoBXH7T26c1gi8IFr+H8sMsDWSNs/QgOL6ttfA4me3Lv3/M5VY7/Co1moIE4SmoMeK9pXC+G/
Xgk9tGT2cU95o5bvvhs48NVyqaIVHT2BS7BFY9ngdDZmO22ooK/mgNjuxn7yuLbvp0dW275ZsfVR
foz+SstkY0510KqfeesYyMv9FElSKtv9xEq8PNRm9AGjdd2PHeskkHN1jNPKpNy/i3jUOL1as59f
rjXQTCeTNIIee3mNSLIVjbMTqn9hIScUK/NLLUqGXTPyBWt+CExyZa29ytWV5y4g3yC78H88Wqn6
OrWVBaO236d19lqhOWpb65hjlvRnnKvJPI+D/XHvPZ/rn2LB8v2U/bbXQfjcHAaOs/dTmMTfUZqt
DjLAXM26KI2f8crXavv75JF9cavn2P4VAYciClzBj4t+2nmShiJQqFav76s50rjKM1RcXSMDL2sB
ygPCCQnl8i099kyCbI06c5kc4h4N4WQJwNnRwsefn3rTyFJxdDTZ/AoCeYgjrJS2+R5FmHQzNQA1
NHe7EguqHJ/Ua/y+Z3xsAJCu0vPCvaTHkZoAUIFgQKDM4VBLcYGOe6CqSvtzPd0kvoMP0cSU/2pe
sVQxqf5MvEoVzzaYSrhrqLZja2SXZxSAUEV8OKfeHCEP5y9ZyzWmRvbtekH7KRQDxVXqsX83nMKu
54znYeNpcZvvAYh8HRLCkVjzg6+AHS06OQupHb1a0WO5PgQIJhxhdU2RnLkcgp+iyt8JjgAJykIH
Ns6MyEGmk2cWN1H15PkX8zNHPFD5MdY6XOZdpp0umm/+eOxpnSs1ruiXS3x1ULmENlYBvvbFdHxE
L06n/M4eHUZqqQmEdZefsssND5sX5RtMNIWQOPzjTEoFkAmUIPlTRPSO2NqM458oBZu8e8ycoX+z
VRTIerpl29Gzdx4znOv5OqsndXsPpy4MHMHBz6WCD+PuJ72isOO28Hpf7iC8Rq5nnm8vGA3DgGtV
+eQDs8i/2mD54UhVut+udRZNa3K3DXRs1vPwaU6m+mycn0f5ebf4HNJxW/lT8e/QkBg7UZiNLt2y
1SZcM2h7F7lf8EXpwgXSobLnWTgt7QEWiop05o/x+SeS5crMQgLhJnSJ0v03PpXDVkM4rVL1EW8J
xD9ACTGHoVLPrm2zHqriemGJjOi6HYh0LeVgiY/QfMFHEaVL3V6y0hc7xJxKorcnv/rjzHddFlgZ
WiaRmakBKsKBmA9H7Zlcz74aQkDU6HYmGF3xyeSoZK7GLxAVjgReppRAa5Eyeg2Z1cRwzibLydMy
UjUVuKGZPthYymH3W/sKZwVxpfSYWrhBcOslHtWVPwNZmPYE9K7Se38YlD6KQ7OjDAnv4iSnQ6sK
BfkrRlS4UdcQglEpDpajhyMDVR1hJPOLM8a3iQQcpCp1sIrUD35t2+9HmZzUYo4wdkFRv4BdCWY+
XRcpfGqNRPw64QACaiCvg84GjByq6q6xJIPIsnlJAeOSaUR/EJ9mR0Bn8/6+cSLnGGX9pq77Sjpi
O/xfONWzM8cipsugbpWpF4FI89iDCcHc4jp0pxQma5la5+OEInetaM7Ity/qOf2zXzQAyAvwf3T9
9IPB1yH7U8q+kUSu2AlB2Rvh11kcZRJkwF7W2P+LwZwlY6lZhlQXeEMhKuICola7l4e4SjtqZcaG
YMtgxOMZ7kHsLoih8Yj7ECTct2v+zb0Q0jjzRePyFj6z/Mc/nYy0cg0tSRDj1Y/YIEfCNoedTCOD
xc7O0d1LEVIZld9YEFBsj2Qi93Nt4SoHrTEtNY492b8Lr1vcPyEfi0akmFW1XvAUScdV6g6NbXUj
XtcWXuTld9k+CzePevRCE7+0MplsA74TZSYtoBxqHZLMJ8oQL4feN+4bcDF9DueV7PbZxt7ZAG9o
4ys/VngjQaxXGTYD0OpPsIjyEn2StXX0QOvVrTeL4ZSyoSUKDwSTkYDZkitBwVlXzoagGI8u/ZbU
Yfpf3VP9HZtQBIpj4vTrQ1aEpiWGPt593tKn066o6kVVqVwrPAiT17kmtYVf7me0sZA2tNT1izon
OHKCXTJBWikZ4dOgN2EwYirhnTL7B+ASImfN8gB7sy6Oin90jpgAFGhEru1cZdT2jlNZVVtKKCRB
N3A+s2e/HZ7juPxf1hIpYQN7XEPrR7Rcsr09K9RZgEIYL03vfZRWddrTB2gTParVJMC040Y2eplp
yNO+kWyWsmExxPNLZupb0QEwNlashJxUa1Ek0ZBJux4QVCF8AU+kmXhI0k1U5bU/bwwJdWq8ckns
ZKaYabEXNRhrCo/KH8vAuQlGG5Z2Prkyrez7lFzBfmLYJljQwde69NTnPmvc7xVOC4DzojETiUvF
yf/lGzrDwruzsGTfJEbkb8ASZ4WNqs0VFSOIW/+KQNscszRdAWaqVua55TdYMU51sm00GhqbV8hX
YohbyN2/+VRlUcSlMiP7I+coQq8Ys5THDj6Vqum9BUE8hloZRhiXlGn0WkrbfYhYvHPCPoBfPSXa
IUIqYs7pGyKDnSw4JpZBlW0gM+Gz9kRrN3Tqp/Nb1Md711yDwrgtHruGT06y6+Nwkqps6jeVT8k8
4fo7BLSykmo9dwCJmwNZxOJLqrcXs7HNlJjSPysuDv4b2aj1ywswu0hZBHMvzLLGDYg/LRiLRfXQ
KoNZhCKwBFQc+pdMUHUMimWfVfiAiYUL0TTfaBMoNwDFci+C7sksXLVzjAKNGIfoJ4ps8cN8bHnE
fEuOCP/axSRcPvgUnnrDzedpfXHh3bJaR+o+v4zNsM2oBes+ASL2pmitCwbAw3uA7EJQwW7YFmCW
6rubPuzy53enuVhokmWbjMwtr83AEPh0WWSmg75CYxTKMSbuUbaRP2tDNCan2T4V7+Saz9/y27Q7
b0SPjRtNh5g9yxAOUlK4qWZ+nKpw1Sj4QkUzJkOzb74XgQ6FBTk8IP60n3TdgZGUIDkBGKXaJpXN
j5Q5Nirp69+XLnbMZ2VGvHXsEYtijujgaLDis+UKQmozVXUmtouO4bKK8lXbY5m2UkdHVaBbPnjf
IpLYs7AgMEtnIEQI6q49CaW3dUfpZ/L7PhKcX3vRWxK44mMs6PLVtRGpmdmgVKyWEZPoVfv0zKWi
QKbVxxs5KvI7d91A6S6D0pZj6hQkjNWooqKXCbQrbqXUTdFJoT6czMrLh6Oxl6LnvPwG+9UKsBPM
9aU++supJfnfJQG3s/8dga8buzV2iBqhbcwmesvmLvAHmBdLjTNdX0rkAKSSnhAnaTIhK89P2Qg9
jtZ6nVtsArSJfg6I0M4dHk6/VAyNN0Oo0lhoU3vOnq17sqPTWNdw8AX7DvBXAeWUYDRXB3aELKv9
tpueMRihHrgBj/uhMpfWUaQT0+MJs6flTYRxXZ0zYgf/Bd9rZ7XUBp7aJaFLuIu43OHSBIwJjqKR
Tf9H3GD5Er8JQEsiijniNlKtA95WYLyIYr6pMLnYcIPPl7vcIbW7ZLtMGcH5H/nIttkMZRWrIwjI
99ar3ofWyKVEFYd4pL1iQaUY3G/e+7+I33HgxaRzeYB7L3ACdXS3GWLbM3JmXkWFVfAMb+xf0Iyh
aD+5+FrHFUIICd2RkixsB8FurHWmV0ZUFji3vp7Bw7RnwSDf7cOx28KsrFpcGt4ozS93sqNaJ95M
3odJCfPWJprWPqX1yvocPdXzD6ZvOPzEXNHwUKZAO9TeqXn+AKYwK3IWBBDJ7sFIvQuT+RQ8wlHc
vipETcjafQm1yu6UA5eOf9ddxV2UGO+MhAadnB3yGtIlFXjA5vG2S4Mq2jaIMx0VpQma36YFhifi
eDjlTpPaoKSQlWlGSdXf/YbDzsBpbVOE5wEjvsMsQswZic86bG5vD3Y7YbD5qiVZBJttALUqbKkL
F47QlaaLVlla+ygkYDZhGEqwj++UL7tKq+Gs67i+b9dk840pM/wBHazW8frTjwhmjZb7kkFT8N9x
T6US+BaLFj4tLxDdvMccTzD26ysENjbAsbQ8EPX8nh46F8zY7AExpDhyjOVjcrccgAxLgu3lV7dG
aHVeH4pkpl2tUtYmv/tH3sqcCpsrMK3Mu5wZQnRsJEO7Rgee0ef+YHrbBOjkZp/QXTH+y/UMtQyy
LKTWnot/UdWQFjQ4ZCr06RAy497bFnc8weJ8PiOWKegMOIdtnbR4M5ftwhsErr6BQUeXykjoQk2x
Ss1ZUjsiGtxEJi3K0MKvWdaFLlaKdhZq2IadPGO9eGji6IPIwZKK0lRth5fnpzH7spxBjiygA8Ha
XI881rQSFDbNHnOHdtoz32bd+6+TOegZ1VhmBxuKDLU9ZT1Ho3Uz6LB4Ov4DWTy/VFMB6YV8uv2V
3ZetuYJad9j1TsXUuMJ8b3NEMeZF9HuvIsHvnSkF0COFw0u3ORldYoQZqFMeqzGlppi78XkNYddG
N9cqLJ7UIcc18S530L4CIir1nUTZFYrSWa5Us/R9kff8pgm49INEMkIrAiBFjnJQ/Up3OE170Ffi
K3/OfO/ZPoBAb7Cc4ytYuOuQith5zpccfRZxdcJGxzEFyBipeqlnVWl9pMKLfaE4cVg5M8PfaBCt
wILqP+RuIKP0X2Ac9lPRWEjUCp3jgrMvidAnJwa5oEWC4M/EUQZIfWD+jbF8qlnZWm+sbO8ffgw/
78mWxYcQvIiqozKrgFWUZt3opgO+1EK2bfpkbZ9VZ9B0bb12sEM+fRcopBYpTqwENhlVdSISraJW
fkBX82lnFILq4/BiWHjqzpHF7Fvc6WrBrRGcrKbtH+bLPLoI/5rUF5t+QquG//tHhprNoPi+itpj
eJs7RxEOWPbiDxW/eM6ulTC0oBd3WlJjxSMuOrAzCaj4vscTYR/YV5Vyg7OZbzWdbiAC/MOw/Sd2
YoflzdJSXaZf6XhFTOO00RsMhmtXk1yyh10bH8LNsNjIn7mqp/s1V3cq9ErEyGZ7G0TRd2Jpgeby
Hbhwlf7qDgtskV5ToQhydppiCHr82LwU0FWny5G5D7o69PSmZY+w9VTIrns6JvnEmBR7kZ7E4wGM
IChco2wfZKVLJ6PsComMeV2URYFzVjfKQmz6IOE+oLvo83SutLt8vfWiMNojjpyhjm1D784e+gGm
prbGACDz3sRph08Wejptx8e1/Xn7ZPFihKhkGtoNsF2/H51nAv5tDcwbYtkYx+3aucXQi7UOWJFr
ODQVbLATq2WWqFz4zSx+w6VUT0umA+5ILye8BkZ5K0o4nS8locxHxr9r/R2ww5NG15O9uDekyaxA
y4fbrBzW9/3JR4vbmdc6MKEI8z4rxsDWG3cTomByzdigG7hYCq5K48n4g2+0L4TdmAfvsGGjQal7
O0x4gRUrqZu4YPWytbzIEMiiqd3fUI1UkJiCqCH48iKe0/NW6D6efcaxqZVbUV0Sr4rJwlBTvdMH
oeJVGJnowIzu6tz4huD8Hi7e+o21TX0g2OOViHC620SZuNpDdzmL2lRCItPIKDYUwZgPAi6uaBcf
+tM1qA21gX16pu5Llr3ZZI1ADR5K80Rxa/IC9MwKriiiwFgZJ/fR9eZto4fWfrAPSjQ6shNjifj9
WY6CUygJOAljsHsFsHykf/uC8urhmhCkSd10MyQrQThcFXqMktXXfOWSM6kpNtWgDx0XXZNV7grV
iLeTXoArVsIpqPwFO3DekUGCIIl7+q7dsa7htEkCZCVv0KDdWXrSJUyyR959GKhs2OpZopUhK5mA
r/D0YxcKUOy5XQqZbljTOroqWNcAJbxEuKZAWS4JY+Y7dBw/Uj/oNkUYxfm3yhvBWrxOHRN50q0v
oflDljqmO7eCPqe8SOn7/aFE9r4A32KkvDNxRTl9/M8JF2iLYrraYbqczkNm5pLN0L3a7Dtgx1cw
ZY/zf45xU+Go4u74SgBiYaOKVNkkm+7ePQKmauQ+4d60SnDVzTZ/EBtNBkTjz1kpePlTLXuxZfxe
G4pGSsUEpAwwPNXf7KUwvy/DnOxD7PzZMBfz8Tn7uhMrw5OxlpnmVIxFtOKI76AVWGsTupR3kIE9
4p9jzI8jFsT/bOQyHdVrgWP7H8cFAmKPrBLiMPRvNxf9EPAvqmU/wm+nI0USQsJAPbcDXMCehdSG
ejci0Af/E3EpnFE8pfreOfCkt1XzuekMMbsFU6OZqUMKZSwz515sNJ2wGbgHUv9mgGPD7X5HcY49
9m8X6UuQWL/8fM4Dc4jyv7WmtLVrDj8eVjukfTxCQWbPA0jVMyeRrg7oKdx3Ge0ScHSNcqS5t8HA
JX62WbTkkZCZuGVdAhV/pVAnQXd7z10OyCiE/WsLvyLz8iwR1AMzd5RumT6iv6wWpAZpHenPlxY5
lCuOc+oS6vWmCEtFjvn3ZpZLbbn1ICHlRBP5x0VqhIoEe/OAMFQ5iZRx2xFn0aBJyFBe3msY4jfj
8gqRx9f0TzjdLIkqMHywizFk/fo3Euvw/en6UZ56WDBXl0O2CBd7ssWctVJ8S8IfTia6K3hX+NIk
uJ4iwKG8JqRV//zjQEtNhHvCQ6zUotRcVtX2gjAmRf/4dU0iM+7qasgXTNp3YXIndi2oVc6+YMH5
koN6UoBpcXcSaZWoH3Iq1cyx+rjh0a8QNjhOKohDYDDJivoxtmwveDPS5b1dEFeDMwqPU4fwDlBp
PCTb5Rh97a04DWznp9H+bk5irqmkS6zaBfkYrdgcx5y5sYgRMxlSxBD4PbeE0HIYLbnDSL8UJ3Gl
J1XOtJeN3pdB/FozD+vdgmVTvEog//QPgAIfa1U2RhfP2ZagAkmAtIxpYN5kMhLyxkWMk6gJ24RC
oOubK1YFWEpJ+bgY6XHRPvlsQfpwc+gxHlg8nJjXsgx2oZhnicY+7wTagzx2fqJXlCPD7oDdxEO9
GQsjq1eeKQ+k/IENP4eKFiP5pdreCQzsFsVUCNAM6gfomDACas/e4ttw9r55qxfo6g/dpSozyTMC
TXzZc1aOJsS83FM6BECXpOINzcd/XNuNetrxg2x0yKax3BAGe91/XhGECLqBzSBePGqahtByI3cC
JNQzspmP6PBChVV2Cm7zYOyEXGJv2hyQfrEMBgJQN5A3+B/B1rvO9cQ9z6hNt87OvUI6Ip6rO83z
tJSvhd6CLJuhkmhwFMmafAIv1D78Et1iCU+zSTqjfbv3ftn8acQ3uj21dJSixJugcVxus0EAV4QQ
FtpQqEcOxGtPKDCOEQVTXkiqmJACZdGpsxvFDRjeuvvCYILaWW+i1olfsJwKotBsKPpS8nSOOgFJ
vUSpzoChduhJcXz58JY6fp2OxsX7vLU2CqxTk6nj684Z5RHEYm9YIpFeGaDAZnyQkP2MD0vgP9r9
Q+ZWCQqiObTzNSkTwcyqEES7c7LxQx01g0Ixga8qmAjLeX3ykGzjDXyuv6KBJqsrxMM1+VmMWlIz
UivDEeXb9Kf0N5qLghglrF4jUolsDv6v2+T8fytLRv8djMHjOBsGWXhYh1w5s1v3dUWPKc8A6GxV
Dnw7Ai0WoWpVJU4hzHJ5L1LXEDnwZ95U6Jo5lAxzExyBG4diZFCcQtpkUTT+8Zdlds2QjTkpi9hM
vgFiF2DBYTWwqoGylavFpbyYeNPsS9Snh93mCwBXtQAp2iNexPXP2UTCR0yDyhgPkWU2lILW1/km
meE5ZmlwT6xpebo7DrP+rYmCwc+yzL6gqdWs93o2A7Pp6gmAxs0boUs7+DoaqiD2y6r7WefocfCb
anH3G1HwfREwewGFAHMM0vPORmEUAeDoGLFkgo0H5xTjp6Bw00C7rysJtukTD/Sm0wkF4Tf8KEPq
c63vw5i1B3lFFOuSMdtOt8PKOLORSYH3Egv/jO4/OHqbHplEHaU6Fzo+XV0EHI0vnXKY5Kzjul/u
pHqjbpZOi98owE9NSR8RTKXQKIOWDabRs34Pz32gZyB7tNGsvgbqinQgbnUlBULvM8+wpeNYVjve
s0J7haW+oYYpcAd1BamvTfVtriYtXA6aKOCCEiP9AMo3xLbEogRrjZYdwo1pCBWifTxFYiSfSBDN
D0LQEth1uUXweSc2CpAxj0Dsj3bZdmf2lSpfOpJ1KEXDKMyu7H9K9MeNs0RkG+39/zE1+g9M/POf
yXtfROVYXRzab1ESTKLENNgOhR5UyigTKC8HEwdc1ZKOXkbxe48VB6KpDr8gTwX8Ca3n5kSZ0Z85
p5C0zloJKpOqJ/Z4+6+J3lYEJFVaae+V5GS8RMBH7KgqZGUkLcqQV+nAqDYv2fU620eUFommXeJv
hsonOn5uDqczZrwoG7iKFaEDkIxZXkvxot0mRfJop4Y5IteL45Anf/OVsxac7jSkTsQNEcxhcdkT
QG89K1hVQWvUSQ1WaQyS+5zoHXQGUPkjk1Su4Vr0WOvGLl8LvKeT01cqNZNGJEDgwYgamcIzgy9U
DHR+7eUSTrC5y/nmuH9tPuL0UZPpOrw1hVJwDNzxW+1dZ3aMjJ3ITiEj/OTPSehrgF8TkwkkgWxQ
cKrHjI9/Qx+aogsE9/EJK7kGP67Em87eZbtNIkWJGk8MhpYOzStVizrwnHR0T4kkRo817Gj8rL7j
OaIC05mlG/k8MucclWe3lwFvyItJKSU+JFU2vd4TZMWmGlR7gWGLZCXlr1yX1sj5eD0cQjS/vQY2
Mg/cXTBNReZUz77uIv6/Le20Xo/fGKnvnJduhkWt/EvN2xjSsR3Zm4NNtJhnU/qXri5GoOc7Z+bN
yQExbYJGz3UfV0PEWvZHAlt2Ih19aTaTEwxi4tzZk/cmErXMRoI9hqSk4em7i2KdJYKBuUeCgqNm
6/3vJsjBNRNPENWkjRe//37qwbb2Vndd9LRvqJpDfSbHAaqIJZY1zJfIyJ9zKSsa2Z9pnPLyc7mR
D7/ldF6bYHrElemVtUG9ahgOmZDio8nnNHke6i/IBeixUdIhuuc5Ps2IeGmXTWkQt2t33MzIpcgv
FClw5e9AIJKZrZ1x0ojyW42Qds6uGIBxY4nR5ZfdDE2RtuiGk48FzTO/1Sw7GHj9urNbuPpkzi5f
2SwtPA86z7fLugWhmBMGL2hDJcFiW4oSnyq+oibJzSrPnCbjFvBQBftyzJi0ewWLwX3Qosmr30GA
JKCR7zl5GwWyK+VyIjIXcuNamPx93p3Uv9WxtwEdw7Vw/0mCnNXvHzbjGxdLCqB4VrWscujryFIb
pzeWjmdZIGebvZWYBQlHI9bDqqsen6mn8v5Pulfg4AYyLYf2sX+3YB4pPcGIv7TrYAe/+boVt8XF
amIXpdpeH0McsDStZYPuSJDNhyPVofF16f9Z7fEAk0mo6nLRnORfbVRGXFCJPDY2NByFW59taCwN
QJuXWDufVfDGSZkcT3sEg8j3gagxypDNtowTdshbqnl1xLoYOPH2ZI1MAtxm+sDJ6XHfyj8Rp9V2
Q3MaZ48HEjFCNvUh011m7UEPVwaY3WaiSK/zXdIYrMfQoz/xTY4e871HOuv1VxOY3tJQhtXj8M9p
iH84Tr2b+ESXhNV4uHeOU2oSiP9qiPv24zLjpM4dUJxcam3cFMuZ9RcaYYAZWh/nFggnVkFme+0M
SZgd3toHOQu5bxWNuxe/BykmNnK99v4b5/8iyiWpR4P0nCTi7v6tpcua6kI04hMk3fJDr8DIO/Ul
GpByUESLTNhAUYYjZtCFAORGODYeQunNyAX+E2BpV21Bscjcyw/4MPBuSHQ3mMkuQCBDZQCZzzhk
SyeTAbRV7Ie++HvYysux7YViJRQC2Yagx0/vNIJEzbhWWSUyCcPXNRrgDP1VpyosUJzcZpfnhX4q
Dokau3M0MulWknRJY+decQlK6GgaUg8D1D1wITawmev70k31NyFD7c7pWR6kzbRN82NtQ5MlNWTc
CAXtuTV+yrzbt8NzTzeWXF2GGUXXIzUhpUZiDnXwx9jA+squLpiPvEQw1K01SiI0YWvNaVo8Hzy/
q+yz14MBUtFAsQl9CAlN2JM3hNJCC6g07XmPQ1Od8LGRYdlM5vK0CuzdCwg0oOwGG2e2eq1IOqVr
uJv3KIhG94bAOEasdO5yV+uUrojgQRjy2egh+lvuupzpjv123byT9LXMxlobFseQJqUWe/OOtIcw
zrOTXUFO5WED1UQDbgAn7ae7RmXAyIxeTRHw6QkxFlyJYzwAiyhf4Cy7kWxkTpontIC8c3ZJLZqn
duts9/rxsVnZnouKxdhH5UTHnNDER9KHQ3TOhpgzikBBTduKxVn1oXKjHRACIDSjLKj5FSNB0pun
HlQvE9QWQdXGRdYIjE2J0+VfphjID+okris3OWcj46J7iVQNpcR7ksdFnEFjT1zqGFCC9JkC1kuh
w1gPcb2M6uATh48BgQhzH3DQRf0cDDM9HX2RnfQPCveerN/mf6UJlyQeNWBRSP2aEBgWwuEPCp55
S+EfSu5HS9faEPeagI/0xIgYiVZouVCC1Vf3MEybF9zm/51ou79pXXKd9EOJEp7QfNl4siK39G2z
CAujQ6J4JAgIWardo1/3uKhbSl2aSujKhxknDR0R7TY1KnGPcp6JTmO7NhJVzAZWaUrO4X5AS1cP
a2WMq+fHE0mOelBemG48ma/rsWUm4YosLUpZvc+SjD/wcq20985OYQpV+hgh+qgL6zKwak93pVnL
xotnu8JGrxLG9wyIuHTEUklgUEuCMnjUYGuDhVmkWb+DNNhnRTuCL6AaKfZX6lyE9zWw2vJnarRJ
Z28uJ9GD0sh+976MTVUYH1dt3GtuGfAf2yvKSeORUaA5kHrU8Lk32+J1L+/0vO5XU+iRcQKief1T
EntkocDHLibIJA5dBCXTDyJDnWEMHIotd7+0SDRv9oO3nvjmBbH30G26FCXpc/PdO+iR4WN/5c7t
nNogUKUlqhJyFNx5mRqf7gnz0w9+w4ZbAXfgehcFou5EPC1PL3ZUlIR1OXj0VaynCdl5HMWdhxGI
AJgTJhP+gIVXXB8H/Rc0CNc2KCLIjsvhgKcV+uNkvSUuCH4Z93Xt/KmYkU1rxlcH49q4/xPJkBBg
sjeTPWMpt+pgsxzsdAm3SgcBxIUazKdwW7aFBWc+Mt9sx+yAXmCHI9JA3PzzAKRU7tv+3yYjiZ+4
61uI/2B1f1hDno+a4B9Lp9YHtx7I7JMrgVFKMaOaRyjZDCG23TAzQVizO5cJ7FyDGexbVHJBxgwh
fRVjqM5hnhhmLfycVVwXgu28dL1OZGUzkMaJZZ/ntOQ/WGghB56cfCeeNZ+oQXicbOfJRVxqS3bw
UPyejMZCTf+lcPtQxm/3Uiba97aGNG08bzRdjCHRA+W58WFyDPIcVZA595905yLrExKJVM3i3dbT
n0n2mtWWQ1N0J6vbVoPD2PNY6/yfuXfp2KmN90AlCQiYVx2uUkuDJ3OrJBERZPfXsG0P2vdJuCX3
jC2dV93odEaFKe8v/z0t4Yp6fEmzNXri2o8v2x6T3YdyI3D1k89IWYiYuyCdwwqZOtZ0i6UOQ11o
w958jq95BDjWuydo/NZbVrIhphUy7OpLcRPLXNQOqqOSnLMW0dRE63PBFrRYwDmTA6DouB2vScrP
kjNdBmhvxhbJfWW7FkC3GY4wcwHNjk1SlbZuQJr4XLO/q3iPnbpqGrWkWX/K0WqthB4o14feThVD
i+zqrbA2/G/RCclaF0y6+hTMApKLe2KSTL0L1PiVq9C8Zp+5su94PQJUso/4hD/eKYsYYTNjgt0K
HOhvCDzRpnUDtnj+wF20GGPpW6tbzJFOXqMwomRLl31j+m6Mc4l/J05W1HMwMsswCsMMZtbJgrc/
zfCYUywZRVP3QbHnstvn9tKnW1EFJVXTh3HUx5VZdASL5n/gzOw4GQtH6Evi6pLADF6ZuVTjaPmm
5yjsNeR83VzfZ4zUgKSJllw/A5SpCZQ7gplF5kaZ7+QWG92+i8e0Unb+KVYGFlc0Durip1QuxFBF
RCX5RDcK4Rnvr72JJTdbc7ti2uDNpJUejGmJw/y39ZMlbUPL/BWGvUWVG3wFDjhM0xgi/16dIkph
VQyJ4N1Fpk6Z+eD/RJgWKOuKWoub2SZyxF2zUq7SKDiIMVIAwBuwrAQ1YkK0ALel3YeSvYF8Z6o+
hNEfji5WQVZi6LJiwqgMQBWT8RCoX/gf5nW8+S5LTvrM7rfz3/6PdTmkSbwULdRCG7K4dmRkysQC
6tyYGoDBg2cnOj0/92O6Klaph9yoFJwBPa32t7vLFJkf2flLqSS7A9vPb8bZZUojTPUynyJN5Ppo
CA4rXSw3qgjbgd2aramwqDkLybHXSa++iwKak8uRj7EKKijK4gGu2MwjG4BA+tcaonXxz4GYM/+T
D1AFz1jpr/RMBTegE2JOAA1IJdQYHDCawSUb6fOUr1VZXS4cglidqtP5x9D/ulZmD94MyGf5Izhq
AD0vELuZZqnuYh4AeVKCAZFt1OwlvLSIyzRixgw3AqPehTjyHFXyQSD/GTAO5jaPmIQ/WQeFvPbm
+9/csa4fF+8bZleAp2jukkxf13vG6weYNhDJjV/1Z/H8GGXiLFgoeoZfpbBS7cNIMczP8MoJQJ/z
Qwa2iOQdQeTdZaoTN5gOXnoKvX6qawwNSOxZwX4ikMs4+KeaaHZBpwVC2LsGBPVPEIL9eQNeZObo
jouVR0WbBlPlwTdBfSozD2CDvGDCLfSKmlG23FThDz3JYjVqN9D1iskHXcTTyLK8oHSM4ip6jqog
pad1IYHes5M3XhJGSnruJynVV1IJAwEchfA6GP8ka2JxlDId7kg5KX5bHDWQULi/b9LjBIRljKdt
PlrBYwTksLOFT0JCukTOlqPxApEnmYxz94ZXJmY4MvbjCnuWm94m2VHANF6mx8QtjL7S8Ll42Pr0
EqjmRlPrR+Rd77m+sTbEceRTt3O0GdV+5GqzZwwGwB4yBcjdLkbsidkLWKzdFRBqSf0tLCoPYzzv
mwK7BcUikt7ZyW7C9sAfnsjsIGGev082RsAm48CwJ9Bg+F0knkzpo8ivQlShazOQoAkuVCWOerv+
HjUoGOY1yHYvVy4gWQBTAEb3glbO8zoIeNIj5m4SS2DZFc/nS71erqG9XLyiIDVl2JfBCrjQlbuo
cvdWFSM7+Ybd1inZDjhJBF4vllPbVHqmqq74H1as49VtNnICR77Du+WfDrWF+SiRAiW6kI7aJOY5
lsMAoMFUhEk+7KJXSn8bWyjGrAfMdLM0i8pxFZ7jQOvSCBveg4w83Rec43hU+hsMpD4hRhCSFvH3
zxmfHnIPTg5ioD2LLyjTU7MxF8/pnlE9ck4yu4vANUctLR3zTw5l2AIzsYX04yQ62DKDCvLqkxf+
iYre9rja4tMNq2LlHpiMXrRegU4HWCe9iJBOeTBx7FPANGTXPIlfkzo7MtuPeAwgmHkZNXFAozwY
HSzfHVSEoA7ua2CXcmFkawrHN3oTVMV/2h4WynM4QLAJarMS5ufe0GSUE487YTBaIGX8qaveMDZz
y9dRRP8E74+54Dko1aYA2UCYHUwfCFWgS7qrv0e993giM6Q2XuFJ54oGUiGcOaJ2L/Uo/ISmLQ4Z
KyrZ0PylOPfpZ5SqU8lBaBXlKcBCsDVWAZo6MVce6bx9+b2Y0fkcdwtr+qNEC01USn3MrJfIOlHP
0wTeoEDQ1eiYghzL65xQa5x77iHxPpHQsb9Dl+f1KYTBSgbKp46kdLRNnbgNT21v4h/s31LiBuyh
MfS/R+6ALeB3b6aF6MjeLLOyTsD0rsZcYFsZNNc8vtkXIrLbMwinkUplvElMYbiUQ7x7umzTw4k8
YbZ7sjDiH7cdAFxp+QWN2rqXNmUeA8Q5FI3qNgKl4btM0B76f3y0PWlIt3VuGQB6H0GDrc3BHuon
dfNnn1DAcQrX85VC3CJtoVnD+F7U1VdjBOvYiIMXQT9zZgMNYd/xHpPJYA3MSpUwajTs9Sw3L91a
hJ2IG04N+5Dt35JwzVYRFsC8Bq12kmFfp4E/VohIEOdesnz1TF2gt0U4Gg643C5O0xqBF2XiFkfP
bsHGPjHTLR0MwZXnzUWqW5u4EMyDhgxl8tAaN4gMbyWNwivkc1+ahNr4Yd0F7TS+XHd8LrWwYRjL
Tli0zDHUmbJkvfO95k7WFJto23AufIDXmq7SN9O5vR+M4i+rfYnNwrbxWA0s71rN/RwzD6+7qgVk
eA4hF4Tl0nio+WK6ayLyiClyK/ZULxTq47AI1mrEC5fFG72bgVucr8X9hin8N41Tgo1E1X9OypwE
cTnMrQyL/c4ZZaM2uH5Ajg+R1sWbDCEc+lhZy2mLD60FyjrACl0OLxI6zPvUcKejUk5gP5AOHAgx
30mpcZpFJHiS/X0+FVBqg8F0Lj9N+hwnXQWiDF6VDHEFPNvNTJ8nWLvZy6hcz99Mlj28G75Omfp+
wDALfGyauEk5sF2UJ1c/Ldc45R9t/cr8PVyT13juoJMCS5u/W84L8tibrG66KKOQzRpj79/Xd77T
N9YI5xIj4/eZMav9mMX+iXGi+FHE+h39E+KLMnAUXRo6V7gqZE7gxQzde+xmdcavGw6aIdQos5vw
MaPG7apCDk44cp+bQKecOdR+GRZzWvyQRN7r2SzrdtNNsmPIo1ZwsQQFARkzrIJbqrrJK6cvvf30
p/stO0bBVciSFe2at83rsqeffHV/yHsehXY5bvovH5Jno3GDLt1mEy0Fla4bErFecPlYk/tKr0ex
nVcTfWxy2Ao/gIht39gSTvqkF9xnZK+AXG+1LM2ZYMmj91CXW1bwpSppRnvvbo8PhYEswZh+8YNi
WbI3QZzVppa71zcbdeW8ybg6x3QpVpXRzUawU+MZ57nCU04Piosx18lDjsqFkLdIFSK0lK8ft1O8
p3w7YwPjSW7lKcjIAs+52exIYsBvwyzCh5UoSlAP1Cy7iffeBKPE11Ji8oVA+ALeLq54t5FMDD6m
1NS5XGlvodk1nYcOGovKJ8w0jGrpBrSZSe95QiKHa0T4WOv/6ohPRcFIN0ISUv6dquOea4ViWPnb
XATamok8wZ7SqirXI7mBfRidx2/+rxpiOu5KO7o5kiqUtbmOOlaNzN7qq9vNjuZWyk4/91tDBmJN
1wST6DF1w/CDsprRtV/TKjldwMh5DOLyiYL7nKSu0OkbTKNPvZ8B5Et4LkmRmaFD2hq+stblZzEQ
EDuFkpeWwBFGekRbGyad2w32SYD2/B1BvB+0V5ZB0Db0YFLz/YxThbRlkf29O2ZpYNIWrmnQDSgt
zi/2bSeKl161c8kXFSb2BYuKpHyCy8riVfRskNJjDq5iFspte1ZXTUOUAweZFjDbs5diaJCnvZue
Jco2C01G/LW1u+MmPSIWuv4qMD7renJ4WeS+OsERMIB5HgplyyT3JOsa+ACMy4jgYNJutPSJ+C3d
rehWURPue7KoYH4wRVF6oYxQ+UuwWBZTckEMLRTmjUBF6zcqgBfWvrWECauEIus5sWctjMePLok+
JAHGxTOf/atE93XVWZxP8EQ2ixzs32uyVRUwegHSBRLb9znHw/HKmbCy9ki5scgrgmqRasTRCIbJ
dzIjIaXhTFdF3HwDM3Gbo/llQaqWsg4TNaKbKRQVqR5c0EzjPIksQomyepGV4Lp3sWZoPxAgJWOL
CXVpaynhYJWiePvA6rqBAFCsdy5YV3pzq98rEwn3BL1ACz644u7Bu4kjwH8s0G8MB/7dMu6rApUS
9T0ndAK2SsjwE00/qJ+TpDWhPqEdrASapBvMf8psBkXUcxibf9HN1qIJs7E3XcPUPwB78i6ykWi+
rB9wnSAGgj+AaOV655U2FsunuqO24mwIYNHyRyIKa4rRKgWN9YyZDwP4IJ2bi79xOcjgncTinz6g
fVWtUkvH2hm8QFVAFa853MLHxMVdH62dDS9QI9uP+xGRZNPmiabzqYQm4MTSTzGpEw0OvqcQNVoO
8lRLrQHonyJepfXsEQlUX4ub5FtHytnD7hG3o54FPc37PYAvI4VgF68DEHoXBqRDAtMsbrsxrDlE
iBqRUs+tgHBrF2YwcQidAZA403Fm+L242drGwXyZYhbqN9Tw/vK8Hm+oSRZ1ZT+4YZ5/+w0sZtzF
V+jaS4qSYspLU4DznMGztl1KzvahC5Vl55VV1Jzi4Pw4kiQ+BwNsu9i2LDKnuA65JypfK2mRuH7F
cRJYcj+WWLxayrmm2KbCMS7dxQvYKm+r3OWMG+bSqic4d1RWnHB3oKA+wBAazyFb4kbgh+bTwipR
EPM/UFQQqfk30yntX1mVL8wOg3vqEwQmc3lxt8jHinqQ3ZKCQ4cAtpk1FnjRVY2Z2e8sT/bFnoBd
Bh/dzlHRnzCVj1Fh24BGo27xY6Ey/WeRWozoWbCLY8l3P+M1DlhmYAc/D/gEQvN9kpwLSWE9Ofs3
cbL3H8kWbpmvvfJOjEHPkC1MeImWi0YQt7PAY25tqfPYzX8BU3f343DGpELINn0WpWgjr0s6vfFC
y7t0En3SVzXav+84tK11U53jsYFjtGnybDjBbpRmUfojh7WMsrQvzDcscxrPZvjFFO0Rs1QmfLfe
JucvmmBEq1MS54R0ZMBDxZDJzMY3HrLhbvgMrj5QkRvpuplfQdaF4N20BkhdxxFLQ0w+0mQexIpj
JDgd8dcPBJ4vNXe87prLPOr5SH59lu7dtnVVW9CzMzOlPbAsEsvLb3JpFBIHh7XCs+AdSmD2fQ4U
Fg3lEpm7Rl458Pwl7YyhrVWuhCyFneHYN1avEv1ARShRjzIsRNNl4RNg1eeB2GZUTsXnrVYb0oKT
h+TZmOxL8Y0sjrOkWJ9RkP4x8VPffQzS5IOwVELIVaVURfZUYh3dSN2BrokXDeuA8IsmW3Z9VZVx
r5bXCIg1sCPuIEt0GGtzKYWONaZOZAtWQt/pcNiIx2+Yrb8c56MCGhicqrkHKfIdCf58jyYThuWm
jdo4zxF7n0ynviVF7nrZ8O3fzoBptAPpM/zal3GeJ2LqunR1l5OxC4yJlf3hmDspMqCZZvpuy7GC
jLF6KHATNeBQW/+9Z/ondaLRk4q9Sz9lPC+s2A7m9yT3ivtzXsgsvQQH9cmVYAFKPLNlVu0WIhTA
Kp2xx18AUa+B2XhRX6tcIyUb0yGu1yPpRFbwYH1fxMSq/6ODxVSuumhFKZ9XC2Hxo35s5fV2L4M0
Fs1QAUzoGcfykkpzyzSuWBwZkcbmRut0Tyz6N9em1g1eZEi9S2wbW8QWbc2Sf6jfvv0oZ1MgYiNg
YMnHOd+TJb4Luo7bw5klCtp8AWJ1+FP6Cnad9F4vs2ve/CkJ701jW0nn7k9l5iO+VEPIpD6S/fAG
aZy2GHTS5pWx/5PXLBwVvvCUm8hYSQRBhy6NmYUbjC9QHOjsYQCxRAIMqb8RjiIDwFRNrNA7zxP4
bdkmpXzYwiT8sh74l/pV5f6x+sZEvfWhXopVoUbhXTMlwKMgGzl58O8C/BN4YGP2LgzOLhp1m76z
zqL31FXEOG3qqtqhuIYUsqVfRzYihZocz2JT3X2NiwfvhjHMKeY9UjfTfVzoIsw5Os5BG5uYgTDe
q7YZHMvEr/7PitLjwf5iB47+XE3TaEvrspkljAyku12b3ov0aHyMx8reUPflVrXmSTYqxl3H2tV5
XRFbh7HBuXmj8ChFzM9qL7kG7lmLvgYRiUb1aLXy3jxbo/J+s70zq8w2As8neQg3v20tveG7e92q
rlUyleos6+yB4TzHKLipf3kwXscdY/2aX1qgVvnlAPFqyfXG46A1SM8DvDhaH7huJCxa/nwGE4gT
X93+W9cpSbcxBsgmNkNPxy6zXgxFWASQ9MmTHqZqcrfbBYAp23R24ncLKM0NHckfXrCp2iUpFmG3
88r2kB2mhkgl+NSr2XyHAmKS0qfnI2ydyQRbiQdtdmy90Q6j9W9tEPpxXllzJGUbzikkrJ7cq7hZ
ca9lwPORWmeonT4GM/ild2u+EptMyR4X44OgnImA1R5sgkdugoEP5fDp2sZrOhfTSR4Du87P6aOu
H0X0it5UJBU0nS4KtxLtcpLFuIbrwmSN3WtBbx5ffs1Bw089PbxVK1rG4TmFnvZaG8axBnMDFQWZ
M5EcEsEwbBCiYtkgXhfYyNTr25ZQ8udsmpPmUt3xvFXNHoDividZ8yUQzGEIt5fvjx/rn+1a7yKY
lkQNMLsj4tSuILFpVNs3LmKlfZlyKXQybghmZEwxwIjD98fb3ev9azn/mMMo6AR81P3M7JxshPij
L0SIEGYf1i1j/NQrq0c2qqqshJpeUqv8M+i0M9BiPnZaRJjHNTqd/ot/INvC7J+SW/oMJurgZAs4
rr4EGj/bO1/J2zTNQmJmbT/NvnOgyvicc0d28QTj1Z0jWetWgN62q6pa09Vl6J95SWzYzJMb3Mhq
7cJz4pMVn8+CBiVlXWvTIxI63J7RYqkI2r+MO8eaKiHrt77FEeiYhSSRek1ab/gOAEOCHx68UtAs
JAMlQLA40BSCmu5m+DMlXLgHcXZvM9GM7+QrXXQn7Vg+sZYmYwyPVLQVQwxnKRVXo4ntQs3ugmQU
9AOy9GBEN1vwtyRPl9IfILbe8HDfzmuk93oLp4kGEpTNyHxdpEx9KussR9i98W1NPhWr19CfkfWu
E4D3StBRjTh8pqbPB/lgSj7R6averHgkhHr5DjZ2JC53Jzzdtf9Lb0Bq2gTd3Sowx/bP7GkrjDIB
X+Sf0BPbXBXeCT/lcqnVRfBYzSjD/bHO6l56UIAQlIxZP95ZU/YE8gtph3fzTyUB3dMfaQd4XLfe
Qcyk7UtMg3I9D1wGVEqJlqv8PCWV+gMla4AdKRWtS9xSbBOu643HqZENKx0/PMCLXcqaBQM3dqPY
S3S5S6Ju9jTvodyHICcFGwawDMI3Cj2v/M3Rr8NAoqTbRroytgiPci50FgaAgOGDHmEpTJf9NRTT
FgooRrXJjuxITOJBR8HmOr27MfDOaKcz8XW2Dde9J1S0nYZA7GfUAGG18qR/H0SF84Ekhz53zEmT
G5tEDmD/5yjGaSCxPf1H8KmPrc3sou8+hq6wHHcPMZWOWr8N5M6sfm54A3M7ReLswYUq5nKwK07E
6gh5cwokyYGIdqNrIgBbDzf+fHSOHWR9bq4yivvTnyxgdM2+/X486so1Nb5En2llm/Mj+vxi7QSu
Wms1Iv4Jzi/6MWgbx5baV0FlI0FMEh2sdt1MR9mNHDHRgPew+Veuag04JxK/AWlJk6K5GIgpY/Sp
wHmEcWjxF9BArabyu3vCvZtnijytFdZBb4ZwOGq8fqcdBcuoJ31HRHudexmkmtS5jynxQkSH6rgX
zUY8Pb51pSKLLf5H1A0qf4nev45B5H4hhHhVCperSRbp8XgJ3sVEVDI3TNfJ5i0nXFdzFkLiklxh
4Jbu6oCS09nuq0Vma8R3ZkygjRKyRbYcQdLn6zBSu1O68quU/9ggnkFg7dOSWf9an5HsV8uHfZlK
5Tc2ITqrRM9mK+Sgr55Jk0xVO73RYPdH4zOaWlfW+QPBs7VqZu5P0z9kFAdJXpR0GvepTTe6mMgu
twHB0mAVF0uXn7pIOZbYeIOWlLX3Qlq7jifKWmHG0oIRJA+zXfm6DNUgwomhIxiNzSacEXU27pfH
Duvzg2N8fs28/18pnOqvIj66/LZnRCUHXsPW2yySNll3yYstk5FgMozhYf4/NEfaEYgHR70FCVI5
qlfC1+FyuuEkX9QGwLkgm9hqlAqmdzfJJ1AWkgclh+goV4Iv+yOIHeg0v/wvbIk+505orD2mBf4k
2PZpEnz+2/UMKVprqSKXqfQHwpvXLltwdUQa/VEluzENNFaYI1O+2zK+bdlQkTFnumvuLn/lWp6N
b2u77ThBXLzS9OpeY2nGlvxJW2IVjbzAFoVLfD7J5zkHI+XAhHavbWhC7gZct5v5eXHMn1v2V5fn
2i8haz/vj7Vm83hEmR9Yr2UHXn18iD0Dkd+ArTNWumkyOKJFCmPaKOxFolYlPjSsrabinWzAIzpn
GHBtgCOY3UusrOrmALWNm1ngWJis12zZikL/Vv4G+lZJ29WuHBa6BTuk4bmIXKN//g0urjJ6k6eG
dab35TlJRLe7zxz5rfkETkrFHAoVPZpXGDwr4SjRyrjMW869k+D15aZ387e3D1K8RtBeATICE3QC
X1ngYM7JjK9ksxWummQBkrtUqRQJbGuDOwHR3StkOc0Yov1+106uHlQoREn6qNJVItUYFncqQaon
XIU3Cm3F/8yhympdvbaF8396TFarkGs+XNLnvtpnd6zY45LO55uI2TVwMl2DGJ1FOpROK+EnB5IC
6/Q4CfeRqAw2b39wU6sjgqn54YjOCgVAjzdJQipg5qEz4QcVtd91QslH7KAEuKfHa//YxOZBsQnm
/dVNfuwtFq942wW0CFSmRKHFLxUpVdr34VzcJvXXclha7fS1ugz/mNqHtQvc8t2GRGIwUcjQGXMm
eWG6NSTkskuPyFNY/4bfTWYfYBvVC9hQPDXTJypKi0JUNUAXV3q5qxIGNWdK/khf/LEkRgttJB3u
1rAlR4iqrie7sVf4PQP9+/padwnNkruRDpajWKIKRFGwPAwVEewGt+APKGhSImweJHQWg37ZveM0
Sx3UeQqn0bvCgX9ndGwng/awWAbt1oHAb3b/0Y8OEH22rXOkRNmw7lVr+DlvC9HyYh0R0XGxpy06
SQxJMlDdy3czYqXvKa0tHK+pSSJUKuUUJPt3xvUFW8t1oWS374BdO4ZVBsh8N6qA92lYEPLEduwQ
tlSJ39cZLtFQp8ixm3Ymk9QfIn4ttb0XvSaiBOUwOMKXZTuDGecGVlT6/d92syj3HqRg/VDG/1NX
Zbp7w6qMM8f0kj6xh5TFTvCzdt6NCze3ORfyhwA5j18YGFPMr9rQce7bR+Yl8AFXFRd7JAFyBRw+
/wQQETnfruLf9OrB0GsL0qJd86fmt5CQBGiUJoL1CePg+8FLlXaqjLezMx+cJv6p9XnPw/ZjMbBC
bh6iFmC/PmKFWezR8gIK1KL7AcqvOVM+sVnsSOcPkHHN/TFf4jHwYGRldNeJbCZyzXK/AdgjvJkz
Dj2QnT20YRzluVZPz0f+h9o4xEsrxYyINx20wxObHdeEHsWaOkdaFJK6y6dGAo1x0zPwyrqkeCbf
+bvHZmUl7AZBn9hL8iWB/tRJcbgO82cv5KP2aGyF3QgBd1asVrdL5jQlFcbTlgdEhlAXs35IhyJr
pAaDvLL02tL2TZNkZKh/khKpZRtPimjZAVDsxfVz8jCFYGlb3HziEbI2MmIaF1+5a/EtKaePwQZ5
hnZ7ytYWhKKBUkejARM4Rj0Aen00ZbCXghkZCDkTTzjOBY2LX+lL9xe3ijUidGe6Fh4Ta/xoRnmc
YpsvbqutEQ9SWrjWkq85Vh4P/+q/MEOIBI4pCXUfdCm+O2HAHhMsfIvGtiraXq7GxmfgNynpSIjQ
VyI6mW4f7liH/wwOA2RF92pLCjruPPs1Bnlo6d6IwQKmzlRQFnxzkuoYztDkoRoZ1WHJpflXTtmC
ztAD5eQfEZh2HaHJyhXoKIlA4ho/Y7kevrriLHWKVh3twbYPMcBQhHIGDv00ixMWb/CPfvZS7C6X
aO63LmI7T3e7eCRJoeUGywAUGcwc477MLnWyVt7lhlR0/X+9oV0On2RpOm0vpo/5XEfnmRgrinUg
5cl8uyGquoLJAxuiNByn+Ky4Pwk7afODQW2N2bkkDPUiN06LR/2skhBowZFEez31deDeTahle/4T
71p0OlqymKtFUzQcZXNJ685xEkyeNwF9GwV1eiDgG6zyJoZWNFRWSFAEnfGkqM5aZ93/D9TTfzpD
rydhukDw6YGL8YXMu+n+6ewzrPTB5wT3mk5A3rgoy06XVYcJPxfFVJRcClWW+5bORm/gwYZHfMP0
BR7Ekr2KVIrVwquuQnhdlnxuPDAhQkJ+pNXyB+YtSGmbcv86r3XgEYiYRjHAuItRp9ds+9jpyrbB
JtNsKjLlIODxjQ3Uhhi/DECwSX8lqt0N45uIcu/Fzkm6k+CiPfQVtU/id4rCglAoTtmYC4mhhMkl
X7HFJXiV2JGKZWFCyXEMZw4KCfCcV0rKivbdOQtkd3O9crcmYrDkuH2QpxRr0zKq4i2QxSTOtXRc
H6CWwRt020Sgg8kUvT5wZds8G6wVjlJ1Br+cT7Go6Ezpi6+8U1zg1NQViUPxV4RrDbKKEZKd6UV8
5/m3hQHnFKRvlF1DGVa71Z715qy1TPJHLc6NISl+QPrCh+D6yC07pLpoWJxCeCpVArhNWJZJtrQo
b1yI85PT3bBtRgDVr4eg40ITGHbLDTeFr9FnN2STzM4W2j85gAVjLvM4cLngxCuim4Us2cyNHRgB
HMTr1PiUzs5aRR7LoVu8FxQPxmYo7rbGUQmtBY0ymU9c+Z/7WVt2yZofDHk9d5bvMRjZa9fTXAqw
dfHIaj1Lr9+5BI3LkTzVCU2AxwQnvkEYN1fAc+Ey++e7SbW5ylHhPAhe+AZLT4XZDVWbS7WoeiSo
yYGnE0oSCPfxNYAIM4v7hIsYD4gbEPxKv59YAjbG3H9db/66iJicBkLUCHOLXrtbjNrLddbPKvmc
v65CcICyhbflv75YxwUv3s9PBKCIx6fCe0xceFQHWQnJwH18FBsTL4pD1/fkibh4yVuIXJoyI1lv
3oMy3Cj86ooL20rrk2iBoYPYtqJY6S7KK5Do+Wc3TkHxqZWyH3InvC0X2fz2rdlHTqs9IoKWmOia
EgYvXaB0Y8FfvuzJuVjIHs5IULK/Ig+uDC3KlIDwdAFOqaTW7Uj3jGE4dHV4JJXCletwggW4U/Hy
SvGq7c0EU2qqUVPJwzfXjkxp5nNxekWaLiR4G5vRj+9BsyO/Br2Q4PXMY6SYslEKFMOJEoYrX+j9
UF9PmfemFre5X0jBTJDe/YMvhu+G3HtxpMlxWEm8IaWhDVx+OB9llnbTo4EgapgV4wNtirQNJ1Kl
uDwnta9PqdjOufqGESI+4G+mWGxmIis/94fHwn0PRYvXmYSg92ptGjjxTJFWg9c+EWa3kWFZQ11v
1QVerxBOiUdIyYNUjg0LJAm5C9Sl/NIKtHTi/iB22tT1mcAgn6FZzoQuiZ0WVb77zLUud4KClNyj
SqSjg/09OXAaLKkX2Og75AagOXfRtU3dgwsG6huejnUGC8pmZ1aR/xYruXOKleVZRkYzbIWAuS1J
UEidWd4XAwe2Wog5aCLhVpyAfH00WEAOwAtyRrhdyQYRFVLqvlTdtzFCnFiQQ0DXosIcBbMYGyxO
QkJMK4MAZJq6yIRaz+hHfK/Sf1HAGN2fcaivjXM58nyXk7dRPQHGc8DoKIhuz2CMLIv2zO+zOmNe
yYllWX9iYqMQoPO4EHpRPIuea9z0HLyk4T3DxQwATD57+BwmN7PBwaKAXzNBKssXejUPGIOPSPT6
pE6un5UWsTrqtogss7UZAkk5Yg60bmy8wcjlE0qfuAWr16FONgzyCk0EX7klVBVQ7blXUNuwVd2e
fvrRLmPGyCugeEQTCUgIri0ReFA+6rAPPH9jdW7GwsEuTLGQjFHcPGT/9sM714OkIY4yjqOo9jnn
BiXrwtSOQOH5rwCEWXJslryjmpeSivNaOiS2cveeb67kZXoRv53y4C/VEkuko7guH66DqYbXSzhL
tcvV4IHoXvwP5aiSkKYEmnqmcASi0EJqbF54XahCJ+sQISHbcr44PsMNUvyet3bEpmLulcTS2agc
qvTlAF0AfBAj1eajaeiT9maAx1H99ahWGrW9iHFlzX0Qm7Nttu3IkXPuGoyg2/tEktFK3+BkduSS
ygFv70+GR73Bw+Mb24am4Q1oXuVxzKSjgfTIF8/mjOfXD1UzY5G4T0crp8m00hWRGpZIe2bZG0J/
N2t7WVMLGM/UV96+JDL7ZNadzDKAKmivRgkNqY1OHR0GgB5wcKXmSkk1j/FigltWxOf+wZWbj+zM
6g0UEOQo08R27L3pSQt8orw0Lx5Ty1j5vTC2AMoe7PtYiFu7u6CK32AwVMKWbTxV5fjwvsAQ4sZx
gt3nEFe8FWgWHgDIQG98i1+fraKp76Wj2/leMHG7MK/d+PDbil1GmWz2pFn9dxGb5iKiAQcV7KxT
mNvUvoFR7OIhgozcohBJdkPopYr39PbynX73AN7bg2w0CAxKdUTLz/lwvZSDGfCC5ulh3xeW2q4O
17u358cE2JUU3QQS4BLnL3mIK47sLhC4q5gjt51On+gJX7Hc6vGyxtT+J+7/JTLxafI/Nr1KlxG3
z2fz3nh2LrDpJRChgp9dgOzEnVd8G0KesppAQEgTpKMBbu7DxeaW3rW1BALET7RM/NiMCjxSW11D
oZw+hP2aOAUHv/kMSz1mDKIoVLvC7YxS4VPLawsCNU6odfnsTuIWNOoem+hHAXHQWjoC5Z/tvQij
s4EoXFtvziBoEY8wCRGxSnfCANiT2HgYAtxWqC7NzrgiFRHxfjzLJBT7T3dyGFygFAsL8qBKvCrm
Tm8HCkOKiWPETbUb9kr6cL4kG1XA+F09xaTIVj6EvZRAdGs+zHiv3Jv5cHx9NXg/mH0Nue7LIx87
OtcEdo9a6YSLFpurchMy49U+4vfT1KI8CI3VlS5Y0DT6KLFIXZrDEuLwA3Gz7vPqo7feLAne8DGh
UJArPysFaV9lKb6BCdbyFmusgfsIysMk1AsmeXa/Oy3SU5u7ltddi96dFZQ0FJiMP4saD7dtekmp
qzfm0Y/ZZgVaff+bYp4hS+6muAhHUr/t8P/SoOD27FO5tuNjFS+lPUZ8GUC1lJkIY2FE7UMKY5DG
MLIXReLi2r2cDQeLieYq0DSkDydDAnCqoBBXHynCUGNf7Jkj1eQrhHUqzuQ3gHsT03a5V6weURXm
vryzzbAPqgyfunCLdT6+wLEG53GCJmpGsL/R8eRtCI9aexIB2k+v3eqTBX/fo9mISFVrvRP4PQvQ
irv9uzXWuqzXCmTtesMb9E6I4S3KROiyNmir0fn/iHh7NN66zociP7Gs3drosCxAu3QZRKDZpZsu
BC2FWh8Ju5ddN5AkjT4vfESYwnrnzX4EbWCdiSsjQrmEKrY0cy2om2d2WBoqCn0VcPDo+eiBHPLT
+aDaEmB/IxABvaWnD4tHVtFbYwlrsAbZC4EYhadleUO9iBEl+wss4q/EpJx8IZuqByAcUsz5exKQ
0SMwozIMwIh69uQJMU3r66gyIx+j8vmwhRly29HvLO4r51UJMg/dEx3cwO22iC+83z7jXdyC7dqD
1c5/wajHuhjoi3V/hAOgAEdGHLeUoGCHXYickj1zzOokKamryWx39oA855XFHtrGCjQIKBRsVlfz
w6wl7aFFl8Rsqz0wTcDK+yO44gTjyn+qh7lJN9tj1gy4fJ3furU7xy2LS7c6GYVxt9Y517+7mXQU
u1sGEDO7LmC6Z4FOijdBBMEvNqn6RPQwYbPJ3g9fvjw+5opnwytLrlgB1mp0Jt3e/zB1zGx95m8h
ng9RS/HEziOyNkJHlXSn+e3IE/CCiCj0vPMaqY+KC+6mPIPW0wW2N4bPi1bMq1VMA/8XiMcHlTom
S32xcSvzj2DP5n6d/OkEQPVj4/Ygh3fCXNshidCWY2rYtXrGIYc5QbWvyRvv0X7hUuUzeQvhckhk
HeIp01b5O4weD6/9bNFu1N+K4VpQxcvS2teW38Ge8HSQzOxLgDGiTUsRkR+tpeK22TdE+MlYW19S
q2Yijm6d/uPrGfp+9SkoM/Bp4fek7YbuMmbc72eqdOJamkkxYI4ufLODra4DmJbBCxC0QyxKR9FS
ASsEO58bUzhB/bXSq6r3tsrV66spkJeccQEgS4gisR269DE9oDbCeX97mLXsfG5zHcQBAZNHtm13
7C8ArX0yi6VnDizo8Bv6nIP4le6bAgnvN3kokF0SpczSZV3BZMCGhN0WaPN77Pw7XVxkdD+ykQpr
IYPeMxbIx9YbXkmouPDWoF/zcNkkAsXnAKIZwvYszVvjH2BhAEIU2BX7T86aZ9S8n0lSwq/7k40a
fs7DonPVSNb56BocyTUW3Ae1ip+0j6U1x01q4QduVMqOwb3GIY+hcWDGZU0dPXhmIArHk8cJFwBY
fhl/Fsr+rOy2aayK2ji2mj06b7D7bbxO0MJ6N0WDsbZUODAKKEK2H9+XulXWL3dgUv8dBkiS8iga
TRJ73OFTxISNaEEdJxuxLjNrGofGecNNX3QZRG01FrgcDYzuOVRNkddCFI96FmwVGxSxCQmpuBBn
IbKopWWDOxXto2mIM91SyV1YqFPSeJsKgqQUvSM3IarKgjwRLeMX/Gbg6no2EV0SxrqJXYGPRTil
3u83clZjjSH8PCYNmjv8p2ac0EzjDAtVy5j+3yZFIFnFoRSdnDBL/1ToVPfgsUM4QVwILmZk7r0T
2zk/bpTwxqBTAojmzKible9nCML1sArGm3LZ/mR2CzHjb09uvOn7SOEni0tihm7WkJSI2kBg+is/
PgEbOwTUnbK8vFLt/QHwOZyOfvvkKBIs7KtFJsBd/cGLDbZKf/GfDJYrexxY8aFyTak3G2Fa2pRu
8H0pcO6s6kW1IKQQ09hrPC3CXD2mBoCNmWCnAmrevor3bLoAOZVnmII/RiFMUXwrCtcPmKlXQYho
8HVnTm0hcMiXczJsAywxH8ypr9r08ibbvreF8n+P+b21aX+qniwvhHQfaKsfIh84PvF6VHrupTwy
GDwRaFh7SCN5yTjavWsQyvXYkEV+Vb8gagRPTV1MyUFMPctq8CR8gUHINsr4GXvTjZpcCe2hR86k
nQ0OafyXTzstk4cwsbwEJBlCHZyioqz8ssN6yuzdRvjGHmsaaon/4cYIeew2NZk6U08ulKDR8YGh
g+U2JMJ4B0cHJOa265OgCmkjHgvDKzSpF3oLL30IugxKx3563EabvWfPjSqCI3VrWuH2l5TqWTYz
QsCAMg6XQd7HD12/lGBBS+/HNvJ0lB35Sfp5lkWk6KU2wmYkf7GHYUrUShQKU8jk/lUgjzUObme1
FAj6+kKkFslue1UzT9dY0y+3+9GBx/MSK3y28KM7tBSgyvGQlVSTS7HD/Gh4iSkfDxoPFc9+DM0N
2lxvtIlm+dNR6PtxX76IgBqE6JMskWUJSrhEQu/bK6OfgU/C+EVcVsqC5Ep90jU29vrb/1dHrgR3
HJ8XIIhH0pDAWrPqUcI2O8vdRhdSI9DSqCYX9hgZe3kSby3M43EE8zGXXV54b+AEuMfLvcfUvEC1
gjzrJrmN7YlKFsQ8UUCczqjL2YMewpj6v6JSxSW41z4SbDvPPbpvUfWBIsG0/r8cazsYWhvEQK09
wDJP4Hyxa1Sjn+/xMNlC/hHYCEaEPq8FaJlZq8tHUwlwzWwABdPjoIvo3MrGtIoTEZuC3Tu7FvOb
jC4E0E2DVz8V087GF8F8FfTlwfUDi4ezFnplo4zBnLbbMelkLqUI/3x3vjjwpQGoVpd/41TnjMhF
ps1hxcdxgSRTJvAdgnpu3j7+7UEH8xQ+bbmInIzHSaRH/nSYB9E45DpHEFIz2DRkAJZ6JMXmkjNZ
QgpDtr4WckQIBIMh5nqmjrCNPGmss4D5B/LCWSdmCD1tv9RkKGeL4/tcs+H0YEUDNsFBYrqzyTGD
os9df3TZZ0aXwCie1UHMH1zMa8x5LlXn1jNIw0v5putnZnCp/ekJJ/Si8iNOo5LGNeGBqKI3pPDd
PQr+yeov2edbQRzbD1Rto5s39naFYI8sLvoDgvHTv/QumtubkTX/8qexa1x7npGueVnnBibhdw9F
8tY6RluUion2VcOecYjz5qMt9wZvsBdnMWAPd4XRNfUDTd72WrQpqW6Lmk1cnF84vDQ2IshX9iz2
HS38QSn5GXs9dFGt5tdx56WLJEkRigwvGwKws1LLBmVvjyu4+tvJAscqrOcu8lCtAPOkApGd1Wiz
xOFExyp2tNTHoL79ayV8veEOgetLLL5+3U5LzXA2z22bTIRPmIfM1U/amMSXMd3ZylJUHAyOIcBu
9IH8pPS3fK9MXR3uf/yrDmEtBGg3fxkeSNDPhVgynGK3my5NRG5to4Mm1TLkhAOl8v5/rPdz0HSL
FJlsAsOL3fEUw6SBOF0NCAsg7QNLstCiTkTZaIs+vN1928c6u1dN7qI12U2LjUT0K3LPnxu8YCj+
a6F9CkLbKZ7MxPpPD91GJUoiz1LSVfLvvattHP1N9wS//fGO062Lr87i0g1RE8TvvBBWlqBIQKc6
78ZhchSgbwWphrGRu4QXkKBfp6VsonhI/zVRHqyZ+asb9nFuAx4JfdNNIPxOlw5UZ9Z46Xgqeg5Y
tLP7mO/re5cLSBf/wAaB+rOJITzxJVo4iy2OS0lGUg/TdROCNX7B8imkx+lVNvsS0CYurnRyVKIi
bNIgLe9T7jL4efj3IZchhgMv+xiU3hFMfVoTZrnTOtedC5IUgWZX3YfaB9TMjIGUNOHvpuB+k7XQ
r9h9zjMUC36HWS9qkWqCLaoVSXDHdSDAC89OJYqBPbpQ0Ruh90HVSOyK/J1NhjalYlxptPFRJGcq
Em6zPaHqdoZBTIvSpBFaAtr4kH0ZUUAyKVHcl9JBIqXxUZ3qN+56nbiIlkFYqVU3O4WxnnWlmW0x
NR0AE9jUbde802P09sBAZPmpWAgxRPAzYxntSYnkvgQ5wqMyVWpDnYy2cUwCMeHmwvEUME6IOmXP
Si1ykuqzwehzlIZiOSQeIduAelftny3RrsVkYLLitHc1kHTrlLRSSxFU/8DBK+JWc5QhxeMimStW
Wb380P57dbLjHUACG6llahx/nFhC6JzfLg5vZYovfyPZPHaaDGLBQvjembDpv1uEdfvAYlOJA8r5
6Oop9NTbaHjmrphMlgTuapB2qtYdi3HwLA7hrMw275HkJ0bdOHha2679UAduWl9Td8O7+EDPDOGK
k2fIfsNYVdBuhE7k0yhyRhKsCCrb7w29ReoEBNggv6vacZiMhuqW5sssSCSYFfFal8qguk0EQ6FH
7typPSLLbFD8n1A+KcYGuX9KGZQsK+pqfjpgaoml76NyxzkrwaNxOKKfUMLEdvyE68Wd+Fb56k8m
YAQH87MMPzccodR9njdk1CnLhZNcrVWMFTcOLAPE1LsSOVtz0ErmiYU2xsbkUT6ebMTqHkKiri3D
SsVdhVGSGEF3Pr21Ki8vcGEKBjgQdiud6fcsSm6qby44GfYkGffGiJJ7u+vm8SK1D0qi4WV9cv0h
zd+R9oSA7TDsfKv59hsI3TOxLBG6BO6fY4n9lhFaod8slkzAaCKF49FI9iqj+558CFBBFXd/W2Lb
BMz+M0IsVVNie6kS0AxdgQkKQbYdTrk/7FFK2tplpEPYw0YhvRdOj/RnwWf7TQcPN1bVrEszfOVs
33F8efiXho6VzR0SEIzo17abMgcNCNJicfyH25jodP0quB9KBGkubX2iXfircgv7M+F/fo6f+Rkn
SkbgnHalk/X/99CCfsNAvISk52ATDV72Pjno4z3T+//PGA0v5KBA3Q+RTXmxxekBgHsOxWTCWl3s
uwWVa/edmbyQsPtL4p6LviE1UZG7snWvQ0eNG3qhvJL6TvkBdSg8eO7/NcnpyHvGrSL2eDEXIz8m
2/kHDuxmHgu9eHHHyzWmtsEuJDRuMijPaKaI3T0++zpXqhnQIB5nalr9btsXtRBIAUfa2enxAp/r
/l8MWgJVcusZLUlLzNNE++pM0TOp39Hk8goC9e1mZTibFw4Qg/oC/0iYMDs8/AA8H77Cme7kH6Jd
8eYccb8gIDovMatg3V+81v4BWLjYeKFmHvJq2fz4LPjavSrtMeCj0AAFscy/JgFgIV/Ia96LIj0u
iLxHdDVX2Iwuvbaltq2gnp8IySZ7hDSrdbWD/k8O2W3vzxZK7A8o8E+s2C7wz1EaZMZFjhHp1lBc
JUEdA+MrMACed3TGP+gw/je/ujl1dG8qW5Zc5vradO0BF72/sUkoHK1SDkLIwSu2PamnxUrAYhfi
PfASUcZesHbLgVVFGZSn6OSRXCtVjgSwb05/QjsApYPE4teAo6Hs3O4JDEiLhdvCtatkJbA6MGjw
JxHdleBAcA6HBMDAQrgaE3sO+/gcvbyQLX46etVLdBtstCeN+tEtBU4kuiKNsG9g5XDtOkNMo07+
3qCOQmyjAchBSGb0UfZ0fDTmhPxyAGdMvQjJJVTu/E9DQzye8Gon+6KXY6CPWVJsvxR4wt3avaNP
yfKsMDG34ovxOnGB0AttUloNLINDP/QXFsChuSdEW/PZvyX8DVknaxQgDoTi33Tytf7yox2nyYdZ
/84jytaLSD8tvKybmBaFKw+Vp4aSBgxUbCawpP6TJyoPZxLJdCWK6iQ8IG7MSs/kTuA/QZ9DBMYc
7JG83z9kkdnbuer6H9bpaIzx0KqEIuN1/MvuvVwbGhiAhmDHUPhUwffa2sHz9/OtGqZJfCaLvZqb
vLewWFcl2yj5orWMQHnk+L5X6Q6pSArggBp4so61cp19xZacf1ntiK/f1q9dvmKOZSte4HnBlrLg
w3Z4DNIvp9KxyGYCyEjgZdkVyv887TcELAkw3I+Nb9C/jrY4WoSqaD1nzytLF3txD6G3f66drjPU
a4tFRfwNNpeiRg4uVhoQLd/uw9CQCLY/ciXm1YwTXqTX1FDK7cz5gEIbvEwEf/5kVPrK8cpAQ2fh
YCeExNXlEV69knolpyMTMDiq46fW4ZZ+p54CLDez8XoJIv4an7hjYNiDpzcUhAKChxmyRG88e0xm
LlPSnzekskg4BVok8TESx2kv7HhafiBCn9nwJvKHzE2uXy36aoZwKB2OEu6q9THgR+19giNRkBj/
3M8yVRzyVoa8qTjRyxtEu/3CJUt1hx5BfbBjXNGkKDw+Bafisapi+0eXfkXv9R4ZqhXNWUwdp4kz
fHhVCr9ex8aVC1a1D/JcfUpeUpxeD3DaNran0YKB6LNnSXhxLC80FWkUqgJWjZAigXDgtbgbwhnF
4LnAH+Vlr+bmHas8uQOdKYT3na/Ni3tIQcrMnMfjhi6MPqW2736WLxz5z0w7mLGjqE3mbzKriqya
Mkfmccmo6xEP4jAfOmW/CltyE+dYHrOllWu9hpbpVIGFF9uLyoMI+tJJjeY7KF0XCjf4RjxDd2td
8Xgeo9iDa2931j9vDMAB1AueazOBUCZk5pfjjpAcCORRGy2LGvqt3hRhku5hc0I9Jp4nkUUDlR7A
l2qrwp0Wiymt5Ozy5eVcM+jADUmTXyHssOVKMvLxJnxNvfuKoFOht5WPJf5NoLSG2Pa2OOqa+ory
YW3fjlUIWx/+3shuFxA2fD8R8At+UWe8zxjjz+bxQrGGettdpTJUzBJT3t7dWaiRu+MeVJczHFWZ
fG55D2flOBw7ZDdX640Wb8psWm+XZ47QJyONmpEi/3Y6qol8S1ZMxhOseJJkxuhKs1KUYYZQnvYO
EVVLBaAaGYg01EAdJHs1bkEpiVg6Nfa9N7uh36ksKps6gS+grz1p2/WthtcbIRZAUFczSrKzWw0R
fHV7tIcy1FwIpvKB4jbfBtddGQHY6bFgMvMNUhXVkil28K6mHYugsDGW/Hx1NPx+ZO/bs96MA4t2
u7tsRqf1Aj3ExvAGbmZIJnM2e3wyIHJSz/fKQk10K8VcI4YELHGgLBKCQxvG//eLm2T3sQzL4WEx
NcAqnFWbqQsSzQj3qxATb8FG8amF3GVCIcoRYALyNGI/EZ1g9LoMz1raHRG++OWtUmpROERqzufJ
AL6eiOrBj+EARowU2P/X4UidKjiVRC1NBIgclYH9J4FVIosqDwBYeKnC6wyVudhexzUGAfrLmVD4
uwkVP0ek+FgCmfu+hNr2NyhFQzyu6jQx2qiGLSWfSwzdKKAlbCRMmrNOrhvF/aZ7QL8V5OKb60j2
7CcMJ+nw3Zck9mqPw/uk4NeFGOlzNYxcTLqAXuWVFDtHM7T/iI/fFXx5FoUmAuGoqZiGa+QLxU1W
RNs89wlzfPYqjEx58sSVpvCisOa08UHPpNjCmFsctmXRkgwiL9sX5LnsTMtCXUnW2tq9l/udBdnb
LqfG2UN2HOIdGWooRgIpBT4U7IpFMjdZRrqZx64RABOxKHtuoS4ean+HFOP8Y9uEb/4QkNBdfdBd
NZL7+wold0Cf0Me70QZ6uHMywrCyqj8+t3MVTGRod1YqRus3YhZIM06iOvuAeNTxL/eVdbrrCu6R
H+CXP65K0rJI/WjlfjXiI4v5jj6MiR5xzE1dXRo4MlozoxDIb1WFz76yWDAZn9swElTmm2v5MObZ
geadD/qXykASyQmYI1i83mqWawMG37usKo/+2wHiS7xYpku/cjgzvyl+i8uJwsc1rN3C4DR/gs/N
uCpbcYLwRsOJgYf5OVwMXJcqjM75+J/doOO9+kxSsJnON9l6HkEOwI843AXxkCbIFvdn4LjVpcgF
aOLMMowb6P7eJaHu1fCJieIp771FzQHSgalwz4/+D5buAsGfXZjtFRv4XTTrVlFjbulmK5BM+eTG
XqIYaew6zrBQ0ge+efnjl+dPZ9Lfk4rTTre2HGNzcWpzCj0gNQiEXbz2XceNt0fmcAZbUU4GXr5i
/2Zgxtx5Qnb174Nfz6tDujH/9KgxbO1WHln20yg6VhQgubLWGvzZOPPb44dMI8oavizHr1q11coS
ooG8jiYDCbs6Xxdrpc+TkAlVtZmSlgtUyVBdtIY2D0rQ5map0nJkquZSPfElKS1pZovC9pEqeww2
rl952dkA1e7JcURbRrIlHxLhnG8pRWVXJkYNWI26PIgHBdSg5VuBuT2N+vmtmdWo2CxRSMj7g9fe
9CNTTMjXKCxJmBaN3ytzJ/x2Ssq08OEeOCtq2fvb7iz4C3fP/81yUNTEkVxjeFPr5FsN8I1onYKz
mqtA/rQ6HtakSxelLjY48H6xWILhgbHponQ2OpT+Y/THk0y9VZfzdJGhF7zeDi6iv/6T+8FXxIjc
vg8om0m6kSmC7/cUj+k22dTaH7F+dYP2R9QFhx4z4UjKW2KYytEJs/R8Imb9rx42AiHn0OoOXs+t
hmnImURAVV4NLu65M0m0Ght8QBKm5Y7Sabq10Ij6bazOgjDYIfDR7iZLX9A6QfQ1XhofmpTvOTCP
OCDwTN9plC8HUFY2R4ay07/ZAKu3kC01t5aCl4HAGdn67iDQYs/N5DzqAr+1ALYrA1+uipNd1j9b
vNrEWQw6x/YqQbwlefcg0WQqyfhTTMpnQLLMkjrNW4nHnAJAttuSjVDSnwWUAVA7OeQj12NFKTiy
XwW8rY3bJhSZi5x6/UK9bwLenFvzQgxtb+tTD31AyKEZ/mk5dRz6VekKiX8d//9RpZ6OeowhClZp
J3sB24MALiqwuNfWM9/eIBsCW88c+qbmk7H+UZm3b+VMBojFppl5S38lMTTQ7CErcyRLaSH29BUy
T46Ik37KsHys0t4B0duGio4uP7ukrotwN/QYp152to9GYptkLh1hs9hV4XCbusWBswOSzq+bFrll
u1Cespea4qUDDIUdT1fhXaVA7rXQdzaKIjkn1iK8InzBk514JT6mn+kMkCIrhX5A1EMZknSNXEjK
8gUTHmlHs1YVMFNBZn7fr8ugQNSKUS85b6EKpRIFdVcaNNPnDhMOVZ3B99Ip+Xb+ZqnG8NIH/Qf2
tIifNSiESPIyOJrybBYVhL/5oWYmrAyHh6AigshSZbGL3iJcwSGjz6O118e6SAIaIsCqGxZNgf+U
PZZYsgCD9v3HGW3DEQur6U5CJtVeQtiWRz+/gMYIPDtcokkTElhE5EIGvP8bL+ykTdQuCX2TesgM
qLUpWf1EMrJg1akv4YgmjUM4jxQyzjzP2L/6YyYYNZucbiXyLmJG0YEETceB/yGdwsq9oTHd5fEm
c1BKcydpaUuTx3jMxlPZf227A4+Vm8/Pb1HbkCA26Utf0wehfbNHOm1pwf74joMeajVUeFvALXT6
/57AxtHRDtXMUEDWKhjIMFofwNTEchoMv+REVASHgdfnXq5/JCqJ98dLvBcVaqBXivWqDba9ywi4
+wms3fmlPSmHfqMPqDwmP3xVqfZh3OXGZsBMzaIwA/B77xpaDCGYfsvs8z3WFCFdtlrt3mZxqjr9
dSo9rT81rrZVBT9QAwVwJ2Zt1CQ0GeCckU1yjr1Y4/PUTPUqYi86YfDjr9ArjS+HXqUrLDQY1wNR
2wI4cTTtHDUQrOKwR7zW0lO0umaeym97w5f6z7RoI884UkabOKc+dijzTkM1HENml1Lcpee4HC6S
9jz+z4YJl5nrJnVv3XgGHngcGjc7EFp9tfbnCsoEFCz5UGGNDKiauwr+fWeg+QBYdLiZSux6VZQp
O+CQ6QhiU+3+Pw81GppHyyKUB8cb+c+/OSkYzStpE9bQEFNUoC4ihlCBmTemITulHAydvn0scnpa
AlAhUwZV3HJfNS9dgLQbSAcwA5TpkM6RKNIltQ+V/tl71HKfOjeRxGsHqx9gGKImf+Lg/98//fIz
jEbPaQH+BHWnj7XiaxWM/4yfeCXclnGmJH13Aw5ghg5dPuqlat5vBPqr6xXFOmb1Y8QLKI9lkPDa
fl0azsBie1nAryLr5uOeywJtgYP7uE5wOG9adqzXMh1di0umrufaSJ8VP1hifGQgPW0MKPr0FAm+
ewqaXTnH1rebfurddo6tLgWUdUUxlKYYV0X7YvhY5ANTVl7dpxZTxfNoLcGHj+yivliLSV8F/6Tq
9Y796Rt/JUflU8zgzHeD2Ug35xOZFmyunSaKyRzIsABBrJOY4oqA8ldmR2DC4/tMSa4m9+A78Ops
7EiggLfWnqvc8Z4PIWmUOdaQKuEt5YTpQlEbn7NrOucSBZArUJRo11bwjvDm5sz92deHiGmgiFti
jvz+FtT/WRgHIEaeZzgbM0awB+iFWNQzKvEuK6zpP+aSJDzmpVMVAri14ItEa5ImAQKGpxfMh1+H
OCq+avPMc9ujTtrYGWwXmLB2U9F8XFJ1WSIUuTxdguB70uFkcsGtyJ18JVCdNGd26IOQ7BtZWuHY
eBFS8xEQdRvRwGZ0MSq2cit7ar6sK+5343GvlmxXg3A4M4Gw9HGqjIGL0PYDGv2pay4hmA1h3GHO
A4XDGHymTPi0OEabKMhQUsCUVRx4lPuP010BhJyJnBeRaafrW1rYLgEnEyRL8+SUR/kLZu6PPuX3
XlYf72CZRCpwEbgTquN3fMVEakNY6zh62hqDjpCt+Tj9XtlJc3l05yeqGT21y11Pj9r4Zm2dyQ4e
kS7PLXUY39X9QRHdT6kj5XzzBwVt7/s4XHjKv3UpKDJa7WEbIQ9ky7hs02713v2JvK1NL0q+Ec2y
UBfBYt9v3AVXLb4QWZA64aYq2p916eC7MKQixBplbIFXc4ZE5B7FnEqihlSTN1Vv511MxpghX+De
4DjxtjAMad2hNFkkD5XTr/0OL+IVFcHr+z02GjpU7p2by+nP5tRxZUulvPaSaMoPu+pOwotm9o8Z
xKJ6e6W5UZGPupnmGtpNdUR9ZvnhfuOWplUo4tmmj7C4YXUYLTDy3Vv+km8VWA1eSM9Uqy+YOuHJ
084m/vqvnT4rEs1Q0P5uzAs0VIDrzByMu88XTlMPjRM+wOL+TCi2jZBV3jxQo/NDIIbnXK6hPJh7
+KsdFMK+xwAtmto+BE+LrreHI8wlMGVzx49NCT2U2pyFgacIenrRaJ3UGsb5GZIdECx5xFQYqbHY
2wYbt7rQiGT+9Sa3WVMfnasPf9M6Y9nu78LGMTjU/28t9R/qK0EpVmbi/drOCPz+s9V1RXWhQipK
HWVEmIgXFVU3OQNuL7kK9BwfXwMn5aIuOUalGI/jHbzBR0ANmva0zmD9HVasyCFwvN7qKWIi2BJZ
6SDUMxR1GY+0NOhFw1NSUveK0XHage3h6yOCX8lX16U2HxZJJk+uLN+S/jct6wmzPsH60AfNueAs
IjDQmMcPUGtfwL/rAjSj6SdVPcpuTszfHwFZsKRBiNkXg8HFor93gFYltD3ug8RCYinthPBvS9ni
SiMxu3wAX4sXT5J0LGxuiXRQIdzhoJTl7QREgXILeC462ecV7UnsP1JbBgpuDrf818I/3uw+OR4p
rYYuXdgxgNubWel1ZMxvDABF5kVPsjfhvIM8GUeHjL6jY5MSrO0RI+w2Q8GsXPnhsuBz4MiabjvT
yBOs55aM7q32UuPeKuV+5f6Rz7AJJmJcXnE1sw4K1yhw6Xd2roFA1QzbnZClwWYvmtZWtOLnSTQX
KTq1CD38YVqyybst5hpJBOY+tmd+iJA9m5GBd3McL1mSXKp7A5OUccDbyRJZ7gXpxdn8xhDHv4Xs
YY3SsGhyNn18eDsCigVr2ikFGn+Vvnd4cqb6wozDtaSun58wnBMX5BHltesKDxIo4FZCBGVpEBae
xkQjlKxhvdP3fsC8apOUJyLm57VxTmlPHkWFAw3rsAFeA1Jt6EfZADmQdZxCQzVgOPAzpf3A26bR
5cy+UWC07aQFLuPGS9dx2w2zbM4mAEddVwVxANn4r7uVSFgjueNRTr3W256JciQ1PU+Y/unFC0OP
UdUvDrowtmfEjxKOUP4kd1XVt0X/N842Nv+2igSxANeZPuyp/A0il0LN1kW4agZWk1fJUE/Ww4C6
2zb5F4knUK/E50ADKz2yowc4QABspBplbq+DgJkx3LJ2/rHyUn0oEqQwfiLhc3j28qozCjIjezS9
i441ydkcmZWCMg34CLeUg2clJTcYTzNXg47G6cxV98lTCX4b7qC0AYgBYqn/Lf35Viz/I1k7OqLt
w56sE343u1g/moW0u5cdMYrUujN+GwAE3B1zE6sQJ5+s47554N47nbnBahZl1zWxw/+88eqM/aw5
0u6RXZ59WI2DG62mxRFDqmWSeOqsqQ62l0BG32AGGlbGWF3Sqk43jlGs8/8amBTAnjTPun6kD9BR
sYnIbMUIweBvwiJvSqgV0e38hL02pgIBXjyatFIpQ5u2Wb0Kj/H9RI0DXeDLf7yvBmACOvp0uMpf
pmMRaUxz8Smzb4xx051ugBxjQG9kX0qTHpSqxNh2wdcUfup90CW3HzAuc+Zul4sNBqbUUZdkRC0s
fyvYVqAOoSXtG/ZqS9dCyKI3tkBUfxLfZu3cI4uGRiOss3P3xFWXqml8GEr/aP8xP6ZHpX8oamiL
GjhgugdLN9yAuN7tVoYyN3U+r4l/gcZA+T0HSHRJv2NQqxELkaBqggrpNFMdFxUPK0SklMzYz29E
DIfag4FoOw4coT2052V5RqQLazv1tpSTy6z0ZSBE/DDR6YiVfXvDUvr9w+3EsaYOQ0RrZsN1AdoD
Sjaitp4PvAu/k7GHl0lwElkvmcrAUfxTdm8ikTdYfvTOKmTT2oE63SUoy1yoPFnC2vzKqk1BmwcM
y3nQIVay5XbP6eXRlRa4bbOZ5jWLJA1jRjh1AQ1r3hjcv00gVIMUJ/SsZI+9FZn+B924nYBTZ1AF
ZK8AJNn157z8XORUzGX55tY3vaWkctCM8y2wUrF5Gkls1Bo0Q6aSRMvy32UqUYM9qQOZhWzwGpUN
0ptVpN0et0tWhDm1EsYY508b9CQrF8x646q4azOTvZPO75E6piSbNcVn4WsIx99NLlnG0zY3McGs
ltPAWJHWyKtdOVxLfXt/TOOtlLBu8c8vBRLEickJ5S5RMIHOngol4OuTNiDb136IeeV7HNjnfRlt
GNbrE7v+4cWZDdKnxqgtcksQjQFxCf+lJzrvTlODlMCyxsGI/F+vdbzooG/3SKhW36Ybg/W7F6kc
T64QnjQxV7mEcctjA1xTEponyyVxn4Uyqy7JqgBEXWEziIqXX0QobndQEMkJOQkOadXWH86V+K50
ttHsnlWJlC7mLelI5XU7KMjzqtwd3zTx4PVGf01Pe7fQU/aSwtz0q6qjOXIHNtGr0vwb57z2MekZ
YvjKW9Da1qME+3XY8ssTx1KH1VC6RydYQP5XwJ/gTltxVhyOt3CwPfuE4oLPVOFV06RSefTqnPPx
8dffh0J9iPD9A/xjIMeWPmdjZqDd8dIqBQKRc1azTqn8YGueAIuiKos/PXa/prYFZGVWQ7tIsWxb
WFBT2gXMGiIJEGHID8ptNinlfGfF+Znu4zTw2NpsFxI0HXhOKe3d1NSRAk+IO9tomL/3iGT8FQGL
9rWbHEFM9STWsYjE5qN+y21YX/3Rc6Cnm6tGuVFJPlL2KYlf9nqvjOyaHBC07JNiXm4px5YibNzp
AvkrAkA6Ab9af/3QBkkfPbJL82kr4mwX9DI5w2Ae1qEsfbqeizBVjo8IB9lWhDe0P7soauG5ViUq
l4iQz42SZXHilx1/UBBAAP1g71CtD/NoEV7fQj0bWwx5vsTjOIKQTjfzTg/6oo3LbFaSlAE/CzPu
nJkyEni0P24wf8EJvQjTE+z+sVJ113gpIyc85vdd28gA1EvzXBmBFZrf9M0gUjBjhT10tEX76R8I
Q/yV891psXuXv3c3qsrTVV7VA+MY2EptucPfCWuqBAq9jrLzaAe9DN0JljCio10ZmvAijO/7HJyR
SCXYlm/pp8BpzCqIrOD2AntDZsuw81ceRbnxQCjks0WcmZ2nN5vIfcptkaWU8xmvcIWZA171VAca
QW54iSgLhyID4zpV00M//7GtBhpU1G4IUeb1i6YQNvpUPbCZqk9EIZyiJqSo3lINJtoSoALbtTKq
4ap3LFPBiiOSmdkqHWyw4N6fSFH/iSV2gWnBMmgSs83etua+r5PdjtOKU6kIUqufbbSvXGIjHLE0
pqfS871OWmMfpJFUlKx6EN3yQ53A69H2jQLyfAH2+pqDEv8UYnpRnyoroOAxOcu7UUZxdNy1dmQd
/PZdF4qsJGNQkH6CCC1dH0N+voEan9cBKkJH7XgB7sgtyiLkr1YLbl1sDrwGADROoCtRmAqIofxR
esai4n4EkHqofaFzrBXs27cI80OY5uuzAHCvlJkQ1r20PKBNfI/rZxjBxqZaxwbbykJAk1sEaX6C
qMQDYXdMq3jk5lirSZ28ZapsJ3ieqnSUgyJQlvjSMZA0XocY2ejhzlyVv6e3Hi7mDO6xa9n3SaNa
YWvnWNb1/TdcHmZI0f9502aBkax7AlyK2BYOA9iY+BSyTSfCAg6L7c4QoHpQaJWtApOA/SrVnfvN
zE6nUGXgPbWUCR5H0yvRd62qXpf6ubyh4pmw4X4DwA76rNNvUuBDF0x46qK+d3wwvfZyMKygZ6cg
faFVSv++Sr8tYhTXDbbZlcW3bF83sMem2yiHZYqcHLjPhDVX315s0ifA76U/PGT79Xc2m386L4h8
Xq8EeSJ/pA75xAqmPzsbPM4JixJJ1XaJjpbvDF92HLSjoksrA+7R+1FJ/9iiwQanoEDFmjhuDdLu
OknfU6l1Q7NCbZrA2uZEjiVzRSieVia3jNSiQvBI00Rv24adAkCvWfqNmfvakWnSY6f5+PiFHg3N
a5OMcGRYh8ZExQBSmM21W4y3iaQhbogUmqWOE/V1eHGlglwwq4t4ulFScXq1PxpLOIvrXyMoxbkY
vkxMqR5UQjRxrvysGdUOWBlkTYQgm6P2oguA2/wUsvY6TXDImLERojVxu/6XyvD3NMTjYcQMIw66
gZSHd1ncztVfaL/2ya0ZQqOoZ+4v/mLvsj2mJV79u/VLQ3JAk9TE2KnxgvcyWdnWcnSjkJf1i0Ps
zMAR+b3SIz2fvuegvGRiHVvmI+dZyh/m2yHjf0sPpSjTH1Pj3KloU2QWwEJ4/599e82XONFT/SL1
6nB7pwPc2HirRzqkSAHHmXmhFp9SHMtOhvqb3DqSvLc6+WxCLQHOtSIfCaZffX5quRNyNxz4kdeL
9U1XXwyhCf9+dvkW0247oCIfe8IUNRFwc8FgebVdGTd+LLZ2izaD22Krl+mgY35LZLLZWjJ7RDMf
AHzG6K/9f5ASn4ZvwrPYdtV+zluz2e6s7lL3/bBv+EZDViQpdmIsmpWQosbMIJIPpkZxrc0A+8pD
XoQ27fKsB9BciYoPS/JlfHR3Y1HaTMBF1HexxUvV6g1mwxHjjke7bGhKGJj3SxFprG223fhXYvxw
QenZTMa/s0daJNvx4MF27inddBUo2vFxKD3cJCf+2UxORTZ9n4wwW8+eLH4/pkd+m7gA/C0ULApy
ks1Ve2wQ6po/rPMt34zhBo9ZwEyw9eVY63boeuXdmAsMnq79qReoM7TjXue09uLljg7iSMqjf8uF
o/0a00MMV45MeRAJUQAUCzzAQPung7ZNcWPY34JQWcqGEdN+S6NQKVJVW3vGULVW62itnyyZZNV3
ZvZZ5zbbfnxg2ccL8LjliKFfGPzoNHNV2Cq5APXxHTT5PnH6KoqK5PapEu/mchGplVRytp9575Sb
s6TWneWUP+GDDrFDoCnXE4E+aT6gZ/HUowxkRvgRC1jvFcC/El4mGJdA9DDJA4Yw8Sy5mfvjpElk
zUYmjg45Vh4+vtLcEoZRIhIKz84vikdXyjjDvlkjo4K1E2PfhO8SY+Cx7OS0mZGAa0gL6AaCrtD9
H8IKLNZmJ4LklPpy7JIwvJNSS5/FJJqkSd0nbAjWels3PtvleGtHGFzYfjEyK1Tx4jXkE3k3XeP9
DDjqMd66Y//pflO+tAH6IEH5FUvFk2XhtA7Ec5gcwJfTnycl1OF4w3jNriwHrDND1w+Rq0DOJ7lt
BNTlvn6mp02Ah/3Ldi7DiTK3JnTmFiQBSWPoiVr50lrlADlpGaVQdB+KAeg21qQx/6qeV2eekJp0
uYdM6mcZmoReFU1uqibcAXShPO0OZZXwca5bXnxefdnss5n23OEp4zvBQYfQQ4S3BQW1MOaC1FQA
oSc0R9YwrPY8SPWz4D8HdPbcd0UU1uEVQbaxXWhdD80PW3bHlm46kA/ZwlJZYpuHPtbnAfHeVKuJ
n8GjiYlh9U7o09r5mR+hJEK852YP8efrzQNFTRGiAWp4GJvr81Ativer+bT+A3UNY5sT09Aq0OPT
bEJR3gzKgxUiVA5XzAzH1Lw4UyDXqDRFtNpuR47VQxBNWVNl5E7gWdEflny0Z2XCTS6UP43qyNWl
6tqUg7sbF91QM9GONZdAb2xCPDBHEznkyDMvDm3FY03vCeEa+h0HAJWJVzwFPjaiJ1xPZSbmouKw
31gGv7tl7WW9mbp/+eXjx4Fu4ioj4koMvbTalNUPLjzYlENHWqPS2/oD1I0dQKohGAn3ijL31wMm
HQAHe/JwYFlCz9N12Vb1ah5mEz8qQ465BdvyLvtwoMiSyNjIYh9pmpbXkDU6JRd4PjQ5UEhBeXqf
aDLFcImopL02GxedKOfkhheLj+tqq0dk8O9EyCDIFqAV6szmNRG2BnXtO7J+5nehATRa3UpGFrjA
t4P++Pvd4xqXJzZ5JHVLNGGsDPZhd6ttWnPdgRewWlP9QHXFGchXv7k7P9e8xJUu8HCpMNHAI1uM
VsqUuQ7y82FGUnVPng+wrKNfj29Tfwmz/UQu1qOF4BeEq2+GtKTsel0SlipzFQFjOmUXXpvzHbCM
MZhcvNbGsioqYZ/tq7iiQobbN2rVhqT4IdhJt0U5OJ2e+VITGwwJLVQf7u+v4qJVA+ZK6Z3T7Yyh
8xb5m53S78iOUDDJyDMEQDYTS+PgGAaZLTibpyOi4PUzdfTpTNfUGXLsj9w/rg4u4chMVVrADxdO
hnsDHrEYs5iWNFyiyzUWCNx8UiWjH8bFs4Js20jAZxL3kHMcktWnTOfe5QUjf6BvXlY2+N1v6Hgk
M0Y7093eLo6Ra/aIVIjFSwe+qGBtKlMhXaJyIlN50EpsDcK/17744vbNY6GnlLy6m6zA3UOQXy2C
8dJTphJNl+9dCEHwf7SqWPPXGBz3gbVhNCBuSDrmkK56ylF/TvXgn66ctPd8Nvby//5fgi62w1Rv
cxZlh1G5wBBc5cZ2mPY2hkb+gDh3VVgfpLeNkbSBv9TX5bACTld+v2t8uZFqr06UGHvvMxsliLJz
qIvDVR2OW7to0Bn37MtPL7NoHmoBaqYKUYl/ecC2Cm52FBIb+JRaedr3wJVyURy9Iav+0M/i2qmX
n3mhdZY2n7+yuyEWvRlQqalAhHxKJ7kZWgOTdr8IFnt72rxc2xWb9SUBH075kLK5CsTrwMl5H7Ey
Ggt92Z1cT1wpHBXgdqGIYJ7wdym/HBk+y0DWnlItvEN6ZzUNr5Kfac7JfKslei01USGeEbWFvoa8
K4lCddQk3CjLEVGQ5bNEYwA3FZhzJehByUdjHW8lSfn5BRzCp2f5BuhMq6cIUw7qDAhPDf46M5kj
Dpy+6WMcS0IWTnzacfqejc42ioiPJTj1RTvFKPPMd+LNGym0iOXfedct0kWypZcdfW9DqApCoaR8
GfP4s0Sz7Vu4jKIWxVpuBdD2KA1W6zFoOW14eDV+Bsxg47Y8VfqGlegsymjHwdca6IdW4LGy1jde
B5CDwurV+EBHRLzyM5Wpw8kemnZn2kY1YUtBMCTH6WqniBFcXTzg5HDVEdeW44PhBb87+K9mNBdY
txqDoVIzk7ECI0Q5R+NEb5ax8hyLUTPI9JQXuELjTbHZ+QqqHqfGn+vPIqABd6f8O98z6DbAbsh9
GGkeZ/v/Y5QyesUBHgUvZ8fLFANHByW/P0d96D1l26AQHslJem68SiXYZYfLWZBs8AiNwrFcDNA8
OsfhePrWhj2uWf+ACd68O94fjEiAPGU8PZ2/HE6t4ltXCPixsUtxQcTF8ivRQqLjZqyoGJjQ3KBr
tTFRiFYywme973Ss2eEd1JidbOg8CqfGspmHVFeqTcUSdbLZM1EmH+qMMxuN0ami+G7WmcF+ppCj
QC5yq5XqFd69WyOetqHy37Kpqb3KvHjce5AIXimpbt0o7MTUzSN59GVAwtlxyAQ+V/LAUrDAs9E0
Y8kadwaGLEZpYElvJRoQmdKo9YKvEASEN4B7NnosMG375ak2+InUkXDO8I1viPo4nV4ugM6DyzWK
YcU1ioQqfI6rzcFl5G8ZJ2w/arBYOkbed2ezQ3NTdyTLCeqzIu8o/yiRLMmrcebdnS+kFQaVtRyt
lh9bxF4rRT7C12e8FaWk29wxdqZ7RlmWGgLOgzBoUSwi/LJaexhcmweYJ3nvMKZg05Ady1guvLGs
1r2iTefWxN5VmjwPzsNEW7BLjR58iuM0Xxi3TfBk91L1GBlp/i3mLCmNiSFSPMRSKwMyJ6DQ5HL2
tm7N8nixus2oO2jRExmXjAxlOFKO0C7XeXt8XY8lQ5f1S9fgTO3lxVwY4YmaN6gQwn72jIi6XCeA
P+q0M3yoY2JbD2PedhINNy1k1pBuRR6EfMatBPECWImdwYuVzWIR0t2TCr9MXqJjFX7E13hnu1m4
qOREcA1Z/PTm+lzscSls/K9ropZ4FQlD3U+ptW0sKSYJsrlFAflEhwQOA9xCquBph2WILwRQ4zF9
0r48b19Zwxqc9bOtyukf7bqzRG++GyODRQmHyi7ciOOKzfyHDAZppYbjW/+gxEPNXHt5EISloR0T
u8sMNin2yqEqMcMF/6XENV88TNFXMN+MdD3hE4zKbrOU0QMLtAqGmod9aYOcwXpO0pOCJMEvsrBj
4m6fYHr95W+yvqM1Ndi/8EKx0CI/bRpT0duuLop94dDqstMZ0RAt2X0KrB0CtxWKiwDbO/9ULyf8
rr/3t7mW0wS0d3yz+1Y0J8NAL1XBpGkRfWhpTFqbuMAD2TlvIrSu62m4bfm3MomEdTZPv1HXWhaK
ktODEsw2izh0uAvMABeNFH4TCdhdyZ6fDeO1S9myHxaRoI5UAij4nk94hJnYQVWPZW6AznFOSH+p
3jORXsRXZbjAb+/5n7u5AIVsAjrjsJXHsKy9nNItRfCUTz/OegP7TvhFHQNLBpx6l8LjxNUPH29U
k9AIND7gtiap+KPSuesisU19Fw6UPgVSeXUOYhauV5mQ/btCy1RtSMnp6RUxK3vsjsyBVw4cw2VL
oaPQSBRMxbAje9DMneeXV9IyRpAhZGBBcAs6ExLc3f2/d76g/kDdimdXmfKNGqq1M631UWy1o88M
IUKMy52FgiW6cSMZfWrCZ1gXUjLUuXm2cgoIf8McYMParIaURrjJgHc+lgnc3tBFutAueZSqXKue
q9zpkuByh57T5RS2rGKHdZ2+TWJzT9c3zj+Uh9V4uaXIQnybLZiTBn9HXyEsjr8ienKNS7xgYpPr
yWj3e/azOs8bqfoAGxMHVZlAOUI3ueDzfOe53253OciKchKHrLDf79EnzsvJrx8omsBGOv+TiRn1
9LbkAAFlXrjBeX0dINZnOnoxhSQKVFaBwaiz0t139nk8AWlZszfPqVuxmxv0v3IIGPl/6ny/CL+E
ICpA3gjw5LIPER51dNVsF79i6GPy3cC7ADXOWlyOczSh/BPMT0bK2AkvedM1/V0m2oZ7EP1lvcmI
GroMbTDNNXgyb3GKQWHhFsJEMTxub/2b/2zTR380ngSivEDRorDZwToc1bawli5jnhhHCElHCK4h
wnFbw7rn7kQmlxR0eI84/x1bku2U/TZydH8z25jgVy5TKyk9BIgc0Xl4Bbf/lQCIvJ3URgW8qBbm
UzijMYkQwrSIs3VG23apEdEpHFYaEJRkpIYrI8VplgDCwhfF0YWvy3MPn3+2GnNxHppCTqDMESNc
C4xu5+kbOr9cPjE9mLQmgrwOT3A9bk7OpIrxqOuz/Q1m15bhV/RasWSARlY+AXqPzAsV4VFodHEq
vHX+b1xytfhTZTAJ7Z2UTdW8wBnGY74Mm7xJEnfKIqUIY5pteL0z3DwKtGtCsOHgQYGw4bloK9+k
THO+aD8hGq7Cdi0UUsBWjMXnu0Xlh76J6BBiu3SW4YAjdke76ggzvPGQpdqlHyHIZSn7GnSejAOI
g7DZonhZkIDpHvZZgbG+PF0gslQxq8Zj0xy989SKyuv6VHeARx7CuLcukASd5l8CsM/tFjXxVl83
J21eEHvReYeZxbhfcvczpYYe/UpANTlxQ6LAGhL1T1fWik4EkPdm3iHff7yRKAzpyD8DOMAAJdog
vU9yJdA8GDxNk9gDnyCNjscZI6SNUt4D2AJ9lpCzITkLuQ1TinOQdUKTShst20tlJU6cUR65hcju
8L/TmTSkgww4vGYRJzv6Dn1xg1nfHu2mY80VVodtgWjL91WNaksSRD/5TFtnvHY05G/FjkiQZU0E
GuGXJTaZaowuBb6l5lDEpRi0qmvcVjrmYEQuRAwZfYI+DmEuJUTcG/MP8lsC8jMmL1yPpuUaVZJ2
7Hu1Ug35rXvLrdJOJVVATvkk9ttiqwsA+e8MX7gmNmQ0e3u5yZXDBe0XaArK7cR1aVV3fbd47USz
75gWv8Zd6s8OCUkJvG/cDk8WCudwfGmwVHp/AaAcmzum0ceVqSM6VDSdNK05kiVSKzvbrsDtxOuK
zo+uMvq7g5S1sibzXhStwzBOZuPzSYgxTKlcLkdOjfAavV5EIUWW6Oe5V+OhwD7L2q+NaQxSptWv
rpvfuuhZcE++XohHe/FE2Fx9V/2j5NzGsd8amoZ3ehIvj+1HFEBWA06YLW08T4/lJGvbdoKijIYx
eHpPT641FrBDhXVhSpA5BkdTEPPg88w+ED6NbluCcbqmWeCRZB40cICxMyB2OHIP31x4pKtyCzOQ
t1NXa1N8H8sXflBYbxozzkpMEX0IHAPTQUMuRDLetYQnITQsdlZ5kpF3CFRxU/4qVNjdwrKMhSXX
LL8pATZJVmQ6q+vMceNP6FpReYCVSI9AARD5U+Dd5SHnkCSpQW/h/IxNCJIYi5njbgukxlCIkAbi
RhOsAS2vB11gPy6VIIxUD6MkNz7H3DLZMaO4BqlonvITJVntnTD89Eq3sTdKh2Uym6XvQYnYgbS6
wmxjOAkYqsjT3c8hScFrcTy1ApRUZMxIDHcvzYjp9y/EgTElMq+R8iaD+ibxp9fkpzqXE0+scSSD
TaDQqUQwBQypfxjNrVw//eRvEgbZpqzWfM+8ZAHLJHqnAO55Fvvh/d/dAs76iXALEekoTSvjth0N
ViV3cPPzVXYSegJwy2+T9pW3EZnv5E3PhRMFjLu/ZC5n79dSXQxodX7fVbuhIn1hzgbWXx1NG3nK
qGosIk3V9v3PO1A8jlC+1f1pTDzsBq4sMpwBNk4d0vomrPCec/hKe6h7JQQa9zxW5YLrKVnkue62
CDwDuIecbP5WzVtENMcI0ADceZHv4N/BgFxJln5cFomr+FcBgMclVa8kqqAbxki63/+Y7gXCZ6Aj
rtTq0qkfM+/at1m43M803WLztxJJFccdoM2kcBLtfTW6lA0QqmVhDXGxFZtVItuXOGhHBBXjmZMX
1O7MfTJWv3CZeTUiTG92SjDhQnrC/CzxUwz1s9ODIqxreb9mnqA+k7jdLEoFbYt31hSZ2GI/6E9c
JT9kVz78AVDRcXIK4C5Dt6n/pd3xwAC4IpIgDIkDrV/6ijlKGBatrfGYhAxLVAfU8VmQkc/y4bO0
HztXEEtE5PimyET0gZDCLGPP1VM7FaeXI23dOtynCsZ03A/8lcyjR9FnfbFfJU4xm8vrVCzRzekO
mkawjhmzBHvRJA2Aj4r3yHboEr02RJyObDp/JFdcJ9L4urX8+cJTlbK/W3kHoe4D7nMcawVUU4vZ
qjekQISsnqIHgoLLjkALZe2aPQGipTQAaXdrO0qeSLDvtt6qYAMr5b0rkXOj/TR6+hwjlrvJXQpR
JgsEQYsoHnPl9Fj52cXkQfzk1Qd5QOs4tZIiiC68eYz4QNaA8BuuCIAHETilKCHKMVhCg7VjX/pO
dPDIiSNl4wrRluZe+767LhoubRWm4E6hz/TSYPHVb+ml6zZgjJDqRxbB00ZuVfmLYgdly+GFJiKC
iRzb2Os2F9JzUmOPkAMWfPrf2gXODQiO9V4X7Mm1ufkDNuTZjGiBV52ikgI0d2I4JOFXMNIuSyO5
f/ThUSl7cEJfhds8X1oip2+N9J4MbWhz6aWJkdMrt7tS2kD5FfAg2cYSApkPRxxi/sW56KT2H9Ry
lG7pSD+Ai/ZTPSn0G008tGe529PO6ZD6gjwF8eRm8teDKWMuLLMAB0zML3FKakO5atYONatKWl8g
Pc4KAVI1yId6cBoI/4fl4Qr8WZH5hjv75BNZ8OwOhw7rE+PJSaMMpudusvC6YSqOx6vBh+R3ECaP
MTiuR5rUEnrdc6C/cRq67wrE7hWGVb1D1SD31yFuRxPnksSvbH5RNaRY5sf0Q8ezMH+dbXGaD+LK
U9uqbkik1Q4hs+Rip0DGOk6nQ94sa0fnlzHw3poK+eXyd0UfHRTA4YIkjb/hJN7taLFGmpPl2BSS
fmYtmFHksRf8b3JD9VkYttIBlIBLy6EfQDapNw0kFmfXxurBNFoTGYTNDgwzlty/tKmCQNXLlhxs
S0bE5puHpRnEhnlz7/MBGOuHcE1UfGLyN3GT4Lx2i4oHAagZTGQg2UlqvbwVDm6yxI6ZJfkYhxXc
QRSAYDCLyhdJO1bWNAta3kn2BcSnZV3kxANi+h32mtaDVLqrQhYqcTMDH4pbBXyPC8e0kkckXAdO
160ZWPL8rzv59hRgxqQrYvhZ25ypd59a8eK/2iQ0NS2GgConfK6O7+kPR1HJojcTo678mU6isp+T
VJYFyjBDVaC2KLC1mlNL6eIYjfB369LMW/ibeGKl/qj2dl1QEwukgHlKHInHwi6IHkN1d08L7a2F
4T0bXh+PTj8g12AxDbRtDasMN/ZJBrETBi+AeKooxvNT05zy72HyU6SE5Ze6Bo1wFOhz6eZnAiss
4vZ+y0neBdrT0mfayUW1QpOniSX1PYyCnOiCQq7HvavEKhDNRJgMe1JLIrPwdOq6vTv+7M5dFUv9
1434N0Q4zK6Fj3z287EXdBDsPIqNlz3SYaEpwDcBnTZfshCexY2GDiwXqQ6uhgIjD4xU54eT/0aN
yzwFwHhw95DiEfoZMLjpJIvQMY5EHo8vEGDpGr13Lfn7xAwZLzlB9h5M5FzXYs8lUN4Bzu5kuRKe
PEsH86K5GboRl1WhySfdVtGOY4IHlksFrJRgDeOQDxH6rRk7r9H10EGfUKZAlEFD4oa8iujcSdXu
okAJ8gEmagHBPe0coM7knSUHHNdg+ggEn3ePeDh6EAh/c88IJjBpRifX7AgwVhsQfk6cnyxfR9wD
5SahpRnQl6fWOj7LcSx5x4USjOF1FAVLqlteEN0W5OHyGNzOhAlolFSjJNnXLKGg9YdeLoARalyV
BolzW8vD6lnGMKAIU9Gtd28xCYLdBpXHjxVRB6CHhkLMwSsOt2GDj8/tnDpdVqiKHPU94E6ZKldJ
U3nEEls4b+YDP5VbbdMWXHte9ZmU/HLpGnDBKmBYA/+B+UHQlPrum2U8q03HJih1hatxMzACnMxd
GvUDtbjPPEl3a6ruMRplDpEb9s5br03ydqqBPSQiCcdzB8cANIM5bbUYvTlJDq5929+IgTKKLzlN
uk+WDKSXvQ8aJfCfNAUdDpS4W7XqZ3JwFH2vB8pDSkFXVfIDPeKWjVKxtob+CaavsP2lT8OIFaqF
xj4VpROJJfOzcPvMbQmW7QO8IgmTTfZ96bdiLt2cH8HrD6M64s3oRaeDjClCQRdFNPGqzpFBFHxR
qCk9ck0hNgR3wV0X1wnSJazqDOpA9TgM4NmPEQQgkRAgJBXRbcBUJrorD1xnDt1lYjqAXAembecV
Vki947ch8n9+jZLM74bPqW7HGoWx24WlfF2EH8ZD3xM74YVHfktOFTjNNWUJGjc1Yc2LHNqajILd
dDhLQjEXnhj1w0P474bQvhSL0Tkn0H90hMW9dbf9eOQnWI2o6s6NYENW7uqmkkP/51VQYT9HD8VO
0iMlnDulx81X5JJH6N97+3tHyNBGRs7WHEVkuR2OowG5B6UXRwecKcTgvrniMHfdSR+0f5ocDFxk
70a6uMH5XX3v15HSQSncMUrZoXG3M2ohl2C8tTyfOk3ZTlkiCWaxRbRXLSOHrQec0WY/k1zSF8lR
f8u7t9iDJI3QDGaSDYmXgxiQCHblzJkIwFaYL+hSBxCGIYRtZ3gXnHo9siSyselepfhKpYwG9IIE
QiEL65RLDXkkf6qsaEeblGlWteBbmdsetC54OwH47THowarZOL3rlBidm+WNAVYa555LpJmLUWrY
dvYlEprdqEv3Aa583ARFzXl1OBhe3AoI/3ugAOG0iVNu8FFdnfNvQBc+zY1HEnH/o6F7jm1RgOnk
Z5E9aTNQEbbWqn52B4H350F3anVF+T+kSBoyUipmYY4HPVVb4FtXJ9AH7NIW3dmkMLezJYOVowI4
xwocP+vC/gl0hFSjH/qundHMYxA79/nXZhSwmee3hJE6VcW3dkgngSnZ4JCUt02Qqmztg24/DCJA
6cUQgl6cdm4TIzPnoJExarEMbQg10O7dxIPVzcqbPddR+KxF0LFzA23XGEKphSuIt8+U+QzClLur
B63qNVU7un5D6n1CrRjslGN8voElWXXpPBTgj9cvhT5oMTdSDf+vkEpRgq2xTcCs0ydbYVR51UTf
5FdCtU4uY2gkcOk6wgUsuqPjKKgiZVjM/H6qtvSGmFFjorVcdNdED8Q2z29Bhkrs+6LgT8ftNzqk
7Tui3qjy9hHCMfUFKywQDKxbL5fqs4ZrZxJFIqHypN6O0eM+SqY+eoHuurNc2tlOZJ8E4HX5GFqx
+nDL2MEmHw5bZpgrEwWO4N2FaldZzsJjY6xwWMfX5Vtl5zvcmv3RJK0JNAnD/8CCz4pFclMHgdRk
27fHnKzmJ7fAzVjN+VuiybviTETzqWt6ral0V90tM5m11Bj2dGXr5C0lNsYrTo+DFZl84B78ku75
31z7npjA2GkTlWPaThGFcKKj2v512TP/ak5FSmC9VnrrmmQWOppk6y2m3lwZOXXzqeZ0EhShCnh3
k/fcQ17eSNZ6Q7NdquJDb5m0iIxOkgbeNoi79GKyI0We5kxdjSNfIhQrngOWCzwGAzQYPZbITYZ4
cP18BwRPDeg8CQ9aPm7od4EW+BFHvIrsLpKy8tCfy9ItB3kiErSmLXQun8kkpswfu2thLqO7rSWr
Sgwx25WwrvmaFnFu2B41S/7xcsAk5eLZHxNrDXe5M8FvmDQO4S5BpWqXBz0/wDeJU0kOYyr8RtqK
WCil9GNbKtVpsw/60Mi19TQuDxbtyEBLMTxE9Gou2uj/utw1n1mf6p1AL1MEOrTcNnuX6FgXw0Wc
DBQM2HVPr21LYt7/G4l1rxvawCPGdQzRXMnfm8i5qwUKdjhMsgM+Bm8EUIyb+oVhQd4K3gBZZ7+T
YGo8ITsGXcCR9R2xXgvI/D382p7obwDtyEgrPwDnV47lOfCyYbqKQQjsttKWIXWCE/85nDighv8a
AimKR/RB2h08LPDMEdCU3sbpto92g4ytf/4V94V9CVUDOEYAlub2y+9og82/uF7L4ruQbnjSLOr8
64Om2moTRVqLhK70A17s3cmkbV0bBpuM18SC2pW+0InvkR0XDUMPScG09CIgKWU10wPbcnG3a52f
uA4ikz2xvxHxOyDXR6JWM3qhW9GtgsYxiwvxOMOu745ns8wigoLqUxKW3+XhxDkuI/9VhLJNgRGQ
NERV0Vllf9lnqr3RXeVcJz3rt5fdzE0SJtugnYJ9yzbTroL+z0Whz0SbZIcVN6qP/ZW1X4dPrJ2n
2ybz8BipJYNCkeIMgj1wiazTEcID6EYB8BEQKSsrC/DRCScIvFva6ZrIS2P6MeH9pVH4jeEO/VlK
+xWbYMqIegQJD91ZrFGUuBG1AGFU8W6ybxfGc1jLyE0Z5Baa/x09KVMUpJx2GJ0DK3Bgh+Z2s6QH
3lHztr1fF+9uo4zNt2q+Skgyb0kVkFxqgewWL6HiWYT4AaWcdGYCTB8EGrcZ4pTxa7Ys3ibWCZH4
ns4njqYGIjQiKmajVyDzMZmLju5sDKuVoAXXGxkoAaWPv0Dlw149fZmdoRxP4PspXmbZKlqq84lE
Oo7d36yfIsARtxRoOsMZz9p/9KPbOEKd8dU5DlMRDhAiRxDtTxd6PFdC/bw2WDEGdCZq6mBvKnWZ
SpGiey3wA8necWHmHWgW5hgHj62hswdNhl6TNfnSYcpOQCinFHw4gvbKgMDhFPBfei8vTjiM2rQc
q7E3d+GyhSLl3jjpTw673va3EVeUMzO9e0AI3mneIduKFsoofTcRhEqRZtDJ8VeBi943JNliCLIq
zl1DCQIuPMJxzlT1joW3ziXzDWWRBhYljuBtt3u1AyLUMByhQDQQiLy/TnHNHxo6GCN3ZQ86KM9l
K+5pp3JS5Ggj94BlHyYNClwz4hNo8wML8JL0k1YimR71tAVRIjLoDFJjbYDr/Xj2u/QFT7np/2qq
gDJkdvoZr3MeZKnvrzdVafeE3BIuVx5FzVutDgOOeH1FWAtXtg+Pq9mVmgtifdq3QM2vTzf2w0A0
3yiXxYo6cemIg0O/nG2HR9pY8NsTJV0tYWIRNHi8uheN7L0YxKpmMWEcKTSfjnRZZWVRZTsad5Uq
XqdrcOyZ1x+VjPc8kBO6TQpb3c5GndzMDjOm4RlmEmkY4gRF5zZJ8xwTZBpG56lbUsqLKu8g/jsW
LTVuylz92vxADTgvmYeDWLrGgHhsEW0XtdpyKxWz5vSGxawyAW8Q+20NVaw7SZ3+Etfuk7eLmmrd
Ou1ckIWkhITtxKWOh0Zwq9JbbyAxG8WhvzptO2rwcJXevlgFXnpGcMkdF3rQ55ZCl7ARnG8BgbfZ
o+vNiK3X/NJ6HhhwKPw0B5rjRRHJV7CWUkrqoIX3eHTflvsoFNgapMASVsJqVzpsuodlYFGdZt0B
7AVFwVl8FVaYOyKGg1PIROtjzh5dKsLBugTKVpiJ7nhDt9H8JwtaJvePe/C3YWOzxNAUO2rruzGz
1cFbEDPtojIVf7SItcnNPAfb0rVg7qyn48vP7NbhgT3gMUbZuE7vWN/+Si+e4jlX/FktiBkCuZKQ
AEXBi32YISDkLDbC5qZUPgLyX2guS9+btyOs6QpasleMRo9yvmj/wy0n5UniHCtU5BfaurpJUS3s
eDA5IQRasmkeBdKsx4yEt0PgOcpwPRmB1d7M3CtPq4kDyC/0h7+8iHtaU+bIND1fjmNb30mbJV9/
oqd4E8prBeBmyBq84g0VpzbeXwAJaQGiNBsuctOYd3yKLHb48rEvE6EJf38JKjLQceDcUiN8kGNy
FDoxZTk9+mFuVlzSpJwhunJayPxlsTVZLVFq9mWwKMNf9TafjNZco5u9YjmIF+1o7wU3VJs9UPFd
C98Fc/BhWll1g0zi8s995jApLrTxVyastDSYsaRW15UgwKFXN45u/wUdVhaoATWGy1f6t91h/5dw
4toqbVgavg+cVwm27X2PnT0zil4JIXYMg5XWIpDUptn0i9f6QYh6r/lrKnEhxo7yZOLXjyTtZQHg
AMdIfIbupQZmzcd/a3VnjaOd7fudIRmKkB53yzLkHTBNexcROCWPOJBRkJaEKmtgvSxpk9+OOV8l
T0pEV1psVkRKhs7rnZ3lKKOT1sidt+bukQCLqQuJc51w5BUfsvUbIZwVffZiIdAUqa3Ve7jfZz+j
PLDZJ8kEVrnJ6jEXI41Y/1vhXz4uL4mU6sj2DGyGizQ3qhItnOGHqDwO3EjACYduKsY2B7k37/oF
L5/8iJGqmjsb0RrRu+qZ27F4jDmZqGuZDNHDffQTlnZPHR6qkrxKF2JcOPLRq7xcdqdpY/Fkia8c
cwEqimOiaErNFr8yRBB7zzo2aIZVFB8saYtqzXtMAqKlBILLF5i5T4TpkxhqXF4siSt2oKduEwGm
rjMQEpJ+E/MP6xjo6M27VTlto/KhQbXZ3UFfEZFch/FgSZhdKmhHI0wKIyMXTFcw470sRWbo5koN
fnvWgrArW6CLB5uJuOxKQeBS5jckZg6XgmukRLSFOOMQPi2BCjBhjAJwwvtodReN/MCCiMS+qQO5
+wKCUaAjAYwdphbC3ln3k9hbhN7iDU0kvrj+THsYuvh2eWMlWXpoZnaII4XJYdZ9Joue6xKUmq5n
SZFWzaTfHJvKOT1YSrPt4AQgCmqRVHL63W0vp/79E5TCOH0ub76pKpRjc6oW0IDxLlET7BbSqYqi
ZazeqEQbDA1UdhAFITYAC9H9Sfwx83Xcr3Cut7M9AC0RwxyGdTtvO90/hVJOVynyKOuVfcqtn4V2
2aq5zbPB4P63C+YbSLIWZzyD+eizkMLHZ+MdrV34tlRJpt8GTL83+Xunv1piW1P17yAhiIKoTmf8
2sApbMRIBTY/FKxHJPsyQdRICwZ+LtpF+TTKAdH7sCT+jrXcTdjVqZUBJizQZdo7/fNESCV+oQvP
kkTjtGBDoAuQyAA3sqDJufyRAx5tgPlciURcdRqBZoK5J0QsD7XdJKa5qNvGzYz/z8S/ZVzTbYeX
dH29UCnLqHHaP3NYhdrR1o+/DuUYVzmj5M5HAVxAKD0aRO10FYTYL2OcFdu1M7B9kkIUpVjBmCbY
Aboiub5l0PAC+e8iFCch+ooRJ9qAqo4RW16BqvW2HV4y6XrsrRnCMx/eLRPxcr21fO4FUfV3d9aK
PJEYBmOrwMmmRKdISbHPZkWBmikYO4KcQwXGxXAmH4MtG3yIVozcgFPPnPsG1tVyQ713lQEOz0fc
sXgEo4XFb+OGXZB52mU9c4L+bYoHFzP7eZB3hAs3dgUfAVi34I8Ev1WWCwyXqjbUxswuL2whQVw0
AZn6/CEok1iqR8Ysxm9AACzZXMJnRbZgx+PG6QEn+QPglTF39zC8EsjGbT7mRYkOtkioQ9O/49SR
9RKT7xgG2HyHOOtKoBkhsGxuhBKTm+X63LuLwugE+64Uu940ZHq7z9+qaNBUXzUYK3sxs7Y3MvTl
BwJ3SfmX4D0uNeP+V/X6VbYMCeERQntNz7UfDskphg3T2zHQDgAllz4WX1OupcxBHQ9PGMpmoWz1
ju5M3bIq7CE8M9o5KJLzVR/F6H/lxZNtCbZP9OdiFrkCgdYzECILx5jnJ9J6v3pnmk6q8v6+flEo
M995eve4GykF6NW+xBYTNqmfgOVrER6Vqz2ed4EEDzvPDff4l3NYbb5gA7fDwU1J8vkloAwIGj/o
ids8JvuZzn1gki7ADjUo/KmUMIHO9HknF6YDKe7NITUOHafVoKIH1OB4SwiPEKz2YCuCa86fn1DG
krjiWiip2sW9lseRAmt6GP0ssjXyjEEhfrsodjEdVLKGd2itFtwg9mRiySZJFfLW0bvzuyst1RUr
/uDdlFGkqjUh+H/ALwKnJyLNnJmLTSOVO6a259siCyKzhikMCUo2NmBx2zES6xJychynFOEfbzNp
D17kpUrDI5JLmXgIAPzyKZhjKvkB+w+zcbQpgNXjsvsmSuxHa+loH8p78vGpexHD83zgLE0az51/
xhc3uaAkRJq5znYt2hnC1sXRduZ79ZvtHkAsNS5JE0V3rwYNbDsKLhbPQSxXccW6+EIu4gRGzbyE
aKZg8bqC1qeeWQXHFaLpDesEjGa4pwwXWBfmuUcTaa1ziRAnlIAxGnXwnOM9toA8D7Nr8lenEya2
M/gPxZ/WswgMw84RBP/JxPEQAkrACb7rgOson/z0E9h4Akv0VQ0T3RDXkVi/HFdTXM5pn+S2Uwds
PxjHXYq1bYLSIomU132SAWw0pntPUTwPZpC8wWWKuivAsmpfN9eCMDuRWxOffkIMdFhgRWtEd5xL
qVYXc7bXDt/KKBfRviAzoMS7c0c4lHFcQAliEBaOXv/RzxWzgjEN5ILEhvGF4ch/w8B/7sf35dt8
zuJnwtwAXLeKVQS+dm/DI/THMDasYv4T3ggrmLjPECDokDGILsIScBaZvFWYUMWIITks8BQ1AIhg
ViXIR5EdeHk+jMSN41IaS6BGEuyJm8Gqh/xBGTey4bDlE2mlywzf0OYJdXrMww7tah6ESe1OzcPL
jT3TjZUXeRoYXNPA0FJbp+AuZDck5Qh651YYOgi52YJ6w87l4gDDV4ykDDFMfgSzTB/LDz7LriI1
44KkPVEGpASQbtZOQUNXZ+QhXwu9ID9HUDez3Ua+sO//nEnQ9LPphlOiECkUL47ksexgJRp6DS9i
CBIPDok4jbfKB2IYwebEuxr8SLHbhLqeIuvgkXugwCOcaxEXoRWxktgOqY5gPLu/jfIQIKaGg/f+
f5nGXQiTv8R3VB8gAoxx6Z6JMhbOf6fSl3fFgOq35rzZyJkfZUMPtonTdoTEX5qTzU0Z1u0j349Z
AW2IJnpJSCoQ0G0q5UkW5kioQJFxK+OmfolW3F9g6SIstF29gRnkLQKPJw6puXTaPObYY2H5DVhV
4JFKaDWUwtA12ty21MMcXgi7pGnzvLEIz4x3EdBSQpOXlMESbOZoPpHhHL7xLNamgrlGo/CBnLZ9
fCk9dBv9hQc3v7hFbdAagOcGT287bBLm6oPnCL0XRbAd64byUUqfy2Io4XI+h0r7+jUTs2yo0Qw0
fUPp4Nbz+6TQpbV3uFcPn28Vqnui2m2LKWY2teTQ2gX6Al1aRa1IAGLjwIE6Ehb67u+7XTfjW45w
9oTWqJFKLKPShCISHT47HGTqHO8z/enLenpmKktlwszOIsFr/inwuImnBgrS+SNCwPF1W/fgJuub
ZpGjoy+2jMphW0uOmY+s2XypMUasV8GTr/SOb3Ex5Ok+Fi98Z/yVkibSVqcG/BODiYSsXLx5p+QT
p359bXfsYwQxguHh0ZQelhxswbq5DOiJgKf6/O2cLMDgY4nArvlU092aYidX89ZCkmX+pfoAyVNP
zHhlyD7v86WI4TGmFLJ8CrXu/fR5dWpr7y/n/RAnaKUgK27nJkoI4iJdBM95ynWXyHYVRud10IZG
splIeBT/OjKTVrbXJI3YVr4CzCLTBJWOE6bSNs5+qIeMzb3qFYETLguRkTv75RqV/w4PBPBq4ce3
9Bgux+JQgBCYlc1ZKtfuKLMxVT78U9QxbEgYd8/cWJjLw0wM9s8ZdfNFxhjV/yk7ru6emsUuj8J3
3MCNHHKVegIKwtjYHeGpHzLyqUWdyw6Y8KTv+HomMOZsS4qU1sHOr4S5HF8iYnqoM/Un6TOaYK0+
tzOWGjrAJgUary/3eKjqRg6oD24QgvlhLqlfVBW95gjthNCKpE0M61Sw0zfxD9wb8yStBxrv/wOB
q3yrkUvtnKv9bZoWHuDzGX6Nns+aKTmjRh8M/Wye80hGXPiubEcSmktJ8MjHSfhGPm+z1T/QqITI
e90IKDUTqytgGGuhsM4ppuxTpWbMPCJ/FSXCUjyPvNR6X7gmqYFJXv/9R55kP9Utqq4Y54QeiT6q
caIOOhqYAy5hW88YpmbU9rlSa4iBeEIObOX8Pwp9weCa+poOxqBw/YrUn+hlTjhOATo95WMXfqrB
ttMyzhwCkK71R7VGX0c7gz5q33u5a1FjDUHH0HH0cVqvyWIXQzPHKJ9qemqFdgpB9UtRVgTp5eOX
2N8rKkZRbZs+ymudJxwfe9Q5QJ7iaExLtUMlofRNrgmRN7o1L5gh+znDhSPf3l1EpofCAbqfcSfu
Fswz5XpXz8Qzfj6WLv7rYMcbDsEc1BStY79cuZWZ8dW5ELKa/uuEPyVl0nUyFCNFAvkct5n/bwKZ
i8nVNvsqqO97/NU+6rDXSx6qaclCZmn6ZSif8fOuNtjghmR1zN3rqitHqjSpy5CnH/01I0971TnF
DQV+61vMJMe/zOKyrsgRQaEGNzA1dyWAaGfoQY/Zzk9vWb6zQ03g5YIdnTNhozbpIgfsjmYZpkV7
2fyxIERqT39xWX968Kv3u45luqJ3NMs1+BFoBZ6f7JYEt2kP764Rphq1Ko/JbYpAmhh3i11CcCAU
W03NEr1EmK3sZns0PwkBvp2v0nwMLziE39HMzPFBbu/rvPxFe6zFaRxcpsg5QqTNBdXhSsdlLJ10
Y/DVo3eoecqHkLbLt+ck8JMLVaPEWcx4BL5odTm/IqiNDBaugkwwQasUZwIqEwU7jymrOxZN4NEn
tT5ZOnQA4rY/cWFAQZMU0SjflA/tSIK/QPznv6G3aaktLvYd29GJzBqD+yLtdoN5UHYsAxSQ+6FI
foYJjxE/4Kipa9ZDHPjf09D9ZZQA1AE2hlzfAXhaPGbP9tuJ0axffCdnPspuuBn4Ky0ckX0hnnDi
tI4fp2kHng7dow84q4v8hhet4e0PcNr/fpxjrjByKG3e/Y9vSUgyMbUhKPmBe32w5JT4Eg/qHrPu
g5ou6foThobYlwFid0/LfA90KbJIGKWOKlzxuT3mRfm8duoEzwB83VmXMNhs7hutDRKcTA9Ff2O5
niEXzKMjFxkndMDaC7imZUhGXBCupL1bJgpsNfY9nm4ObreQ0XGyvk05EaViw0ITbCgq0UlLMChe
6tbtCRZX3vH7lwL9f5UcwlT0SuzyVHYY1zmMk9/5OJ82qSqLZs9Rlrx7d7nh2ChCLX7vM5ubfYiB
UQVMmXiKOqtNeypQlsd2oXPPDahXTJ2tuUeWo3k/tPURfBMOv7ueMSUn+g09nMPwCzsFfgY7nL+p
PT+kErnewPJLAqTt87l7IPQP0/XvJpidk3PVghJWYBUlFkHStREEvoNnZ9g1YG4MIuD0qrx+FD4G
GCNwQTB2kcOELeFXdfPcxw9EZvWkniyRdIoCoygGMMkIM1/D/eb5jhjfw8N4x8mL3ifChAEfhmUl
CS7NbhlQ9VVwn0hjJDDrO0IoB4iWR0R4vRZecAUnrnySQ6gNtc9MgL2gGW2f5ETX+D9W2rZSObq/
oi0f5HFCXGtE/HqDQSHTggN22SCD+afbT2HJNiKOUSa/+ah+TJvVX/4xj1S8bCPZyk9+c5GaKOnN
K3HJDDoejMPBgrkhLlVOH5UZHxNueFNqgq8lRejQY4V2H+UaVCEBGggO4pNc6o8kJ8TtDsHdRx2b
8cOo907Uv6gIz3U/3GwVBS9JR2GyYshL2IwSgPPo6MtePburr5bB9YSxBSLo+ahle5QXZN8OaSW8
SJu6tMwgNkoB5JNgSxCaBst8zQVYXiaOMTlPtSRSsNcsZ+mfd1sxIaMK9mEUosVujE5jsnGOKHC+
Eq+FK5JtJ1AiXdAfzcbdsQhsEYt/UCqDkWtCTt4wTnBBja8dHcTg0HHTEWciEZq7SFfJa4CZIz0R
muzAa2ZRRyc3Cb0+/THu4MIqHRwl9MM+JAEJpm3hEkzY3ZR1DpTYV6A4CQfz2/c25b4uv5eO7iPI
elMRQRQaWoynq2H1to3m+gDqPWu9D0SUEa4wITkI3MqSQpFheh4KXCG/bVTq05iNpGwxCh8u2R9/
mqTKor0lZC+LencHBpvN8om1JYXuVcqfvHlbYqNhBaOO4/HD1Z0VxjG4wXT+VVE0iNowUHWcdxT9
VgEhAFwQt9lg1LxQOxQaOPlQD/bFUc+C7+P0SuVE3Lr9xV4+COcSRpif96Cg9orDcMrH+NueNCnD
vjXj9ret/hPSqkf8nNxiVIp94fh+3ervO0YIthCdCRT9kyE2GIhIb/z+F90c/AVRC5adBXm/7HOJ
2RRuyDCJSLogPY2Uwogk0w5bB4dixsOjYIq4PJo3i/ow6QAaprmFD1q371xYbfp0dD003I9auoPr
RvJbJvBrwf0G0yQpRYpC3nSGKSG/EtX1hWVj7P8zBiYWcuazsj2nwRF5q01oz6AmlOJVorwcr06x
oAtOJOWn91hAUBsAEK5Pr3FHGXnIeGbpqKQvEB7+C/uX7jHZ7FshbVjXmo/fIpveagpE15UU+3Cj
uWyvgF2xZnGLiITRcwpwcNwVCDpBe2a17AAoKxUD4t3kAFN0ldfQWR586JDRn16mZx+nVwoAo4WZ
Ho/p+sC1Jw8KA6D733fTxddR70hnoG5qzB8mOptDEk94RS6xzNo6azs4oMsQ7zqh2tFfTUxVpzF0
d+XSFDtTEskBnGK+wBfeAPEFYiOVzostv4P6SNligeyzT82sVBfq/5MlXgEufcnG8f3AauCpHE58
vJNbjb9FSYpGKzUXLmV3hDpYV8LuTrrHulHUnjRchEzpk8BGq6Kx1+Pg8bxodrcg1b91YnIxsxoB
V+JOTbx77XZbedcjWa6KKgBK2hL9bdXA+W954cdIivPsmQnXqScZz1PDvF0kl2Jw+0Ko+PYSMYvZ
DBxsl9X721nRSGVoMNcJmHEbCeZjf23XJ2+mLUSZFHj6USz9goR49yXvJ9FpZfLAzxFgG69irnQB
/b/+uIH6OZxVh911GVsexeM92F6M3QWmiNhv2sIOaL/PqIbPLrEabkRlj01enC9Dyey6qTEqPtRk
lOwBfWvP90A5Y7w077D0ZjmUPQU9SYgzS1itlWCjq8VSly/Z9UEjci2YenhKh8XlQoofgDIZf540
Zi5H5q1P+kjGtvQbOOauzf9XQpPMD4B76mc6WuC8Sw+D1UCFrmnziYHaJzGyPm4moEGkDI6d96a6
QPrEdgV6USgy7hFfP1ybc2TzFGaWiJDtiE1T8dH2vpq+usPm52YybSofG6pAh6ycptqtjqL5kYwO
hrCBFMSbZ8m1qMA+1B/lg7HPdpNqPq0W5RL+T1U+RSaAftt9AJsAikfax02wj5i84IdAEFmDP/o+
DbvGd6/E8EnPJ3tBie60QToDMg2H/e8sOp2Hy7Bb/1+S65TPMWZlyurmBo1QrLQbsngxhjm7d+Ix
ropytidniafOPb0yTonPP+ekiOBCbEPWu7xdD1Fj4iDsCAEXr4F7O3N/PULZ4zb9GrWa1bS/pco4
skDw9oz5jsD81Lez46jfitp2/6nWKuZefU05mXIIa7Dm1oopaVZI7bgP4WPIrHijwGbp7v2/HQ6f
3PI81mWQYS5wjrJONtp3ZKOC4CcYrnkEcOMAQBl3UP4qGApnyTVrG9pXEwMRFtX0WZAj9sXullCC
V5R9Y6q0LdlC3/S8r0WbeIgyGFZwCphP+JE6ZT9lRFUINOrnH+Uit3HgryVbdTxPwlD9MtBV+y3j
zkdbNvJm4RyYIHwDxzVMz6Po/QJa/uy0RtxWimBQ+xptRjdS7vJb9OVlw/6VHg2Z5mKc4ijW4DV9
YThDmpg4tPFHrGf/wzYG4/Eyp05oofxCJlZaInnrX8dvUSLKn4tw7lTmdEW3OyPMRYUcbw1MAA3Z
ZXltxBXXczIyhrSLsZ3cUxK5kpP4zkTr5n2Ewn61gDcR7pa1/mA7zuZQD/qpyXoWm8rW8MBPsC5V
D+X2NHbDLEAl7+BBosR2P+fxsM5TFA8fGBFXJV3NrBmTzOoGMH86t9AxfRp88nUEVfr1VNgPt30j
9HP1xWFYLVnPS21P7og1AJopsN48N8XClpSsEJ46JT2aKeVhLCKR9vPlGG+2we+GLc9DDTFHoflZ
GbRpOYlJnuomKukbDem17UfN3RdD2bLoJHuTP+/MySJPRAB6NOSaNFlR3vCsVZSrs8B4ah3VT6Bm
ikWvAeBrRJXu1+x8Rxl91hqMAIsFn3yU+ToZ3cszhTpV4doZYnMwvXQLzDngkjtryNvWvt8dJALw
QazuT5mVUVUQ3akZtFYYcwpsc11dMDLuezo5iD3r0h2vLu+GG3Do3r/8di13PXHE97OZ1ereTQYG
hxbdKfUI931/V2JBajyENBQsrjPc8BfVFeqzySvI0n/EQPsZR4S+HqHfHrmSUupkNFGOAz9Y9DBQ
ec0hTFEDrdVxUYs1OKXgSjC4moNdw09qT3dmiLtAa9/DMNH4Z0m55y+JCSPgZEM09jk0X0pzTx/C
SqzuWWrxtYRa/gPKYiCtQG98//wRWglDJGO8BqnpzLvxGPyUgc5svUuWHI8067Op7riUPhpgzPld
E8g6oHc3nFowVeu80ehzvgNvMpz3ZMTvlvkBF95DXRywZ2GKMs+WT79a2svEG0viXEqKl/V1/9/I
sXn+2KFUb3sdR8XiOA8MWtVfoJzlcxzgtw9YkigL+5u0vrx/rqlqRHe8Zb8CgZMPc1zethSR+Wjb
zG4300xrnX8uO9njFRpiL0G8c77XPX4lOFyxkY1NphSyxazCB7HMyShdV3OVyHjYULRDyI+KoGLM
pSpUwRAjx1rbNLTp/AgKqWQHCXSq2BfZ3TEJjwVQeYmyT3uo/XwwcGw0IqpwPz9ijw5eHdz4yt8C
JTpe4V2QZErwdnOqFqq78yWmVDuBrGhpkpkgitafAsoOnI+bMhdg9z/t6wAho/wWtHRRKvb3NkGC
N9IMCLgJzkWIAOZzahXB/WxUzoXAzUx3tAtGT/jWBLCYyZ5mOm8fR2rz0pavzHEr4LVo5pi98u0V
apxXcKaJkinVesW8taWaf1QCvh1jX3hFvuCmXe7I9VCwnlhdLz9PRG0hGzvMwxMuFFQx3ppEJ7bu
l4N0TY8srWweAzP9vq8K1UdjjIP/6jbuLLTJ06pCJsUSNpS1v6NJSdtHKAC8/F6av44Vx+19P7aM
9U/DcVreOnhLE4QYAoIqzCep4USO1HQfHiIcIHhubGcljEwB7nzlWZb+yAHGTecW/PQ9Ujalg/1Y
SH220tKL9n+jPV/JVnJaCD4r8HkbAnAuGq/67FrRkEMc2j6treb9ZOKUVdvvO8+6m+LIn+IhP+4H
OjQ0u1Sj2eJ+i4rA85n/L0FNGufqTVSo+EbUEqx0+yByLRT69k+W1cSHEhBNHZigQlqCH4OVLnoj
irroTvBex24JhIXh1+gMNVrWeq2i13z5SBASCDHh3XRtJWE/ppoAOSbYwOeRiwDDhSjuThlz+LZ2
4SqwZOWcYVLVngY6xSFESt492CkIezKmlimADpg+H6dl8kPXu/H44V48dn3Zk45kGgMmnW2W6Zrx
fd9748TIfeqCf1XI8OTpJhhsmbq+wmL3mdtDMScyIFZpf0EyuURe6kbl1Ku3BLPh8Kn4/xcB+vkL
acLGZ1Zv0e/p+nOjbKJhFMLdhcYZxLtmGATMfv/6K7EhLuqrTHAyui2OyTV+nmku5hNRp+XoIMZ/
YMe68s7kCFjdefcJ+hVL22jNCN6tJniKvpAurVE/spJmNB1WQKuoxBQrvt9QaCa+zwIKTznlm/oK
m3tmUSC+Ywy528f23Qvd7kQB0MaQ14KTPlcGCR3rZ5mo1IMV/iuj0biuVEDgMO4oYdj5FFlNrFr1
42lWYFzVTxJeLJ8+Gd1SaiNb1kxBtF/nqkw+J5WUw6TDI1AHyKRJC/4FEJ4i2vJXL8+oMIm1e5fj
HeHLBjlT6sANDkCQwi3Cy9rOo0lKS9xEuSvvVUZLELSE30N5iC7g77X6V8xdmpKZMOeeb8ag8rz1
S9eqUhhc0d0IKjMlOkWTvHNlZHh7Xle1U6lX5i63MCFxx3lQZYu/x79S9d1+1VCoutCO/H+fHg5k
0rPn53f4z0PcGkrH+WmdQgXxo0paQ3CUf3ng42lfftGb7hB6SZ24iePi7COn63IpZAo8/lLRM/n/
1+GUUqcuRVuDEQYsZjVW8LERLLRs/bhcX5r+HTieKkWyEpsMiyp+9u9bnzolhl1Wniw2RO/xepds
t6aDzDwVkV9bHtqMVLVkmbmZAeUWd/VFgtDq+oZBAMNi65t71SDEX+iIpFx2p0siwzSbGp9AqWBi
T5trCnveBfDO4p07YbLhS1d0w9yuLQ9zSiqX9U46apeb7d/s6JBj5o8TbKTA6xehMVQgfYjaO/Dr
8FC/6+IGGZrtDsXfUAfToClTuYj5woTwV15Jr6XX/cKEdIJq6rjFzUW5cUOX2V4Go/nfgn+P0EBw
UJ06n5AKpSmhEdugRwV6EAzvVUmR6/MQG1Kr0kj0Sz9ARZKG8vs3IWfrDCOGinUXZYlrfV/ayoJ4
COxBB5o8OzQdOcDIETefMdATJMsCY5VZbU7rYl4VzAtyAsMxZfjOfd8hP0o8N1Q4Wgiq22D3oRyr
bJ40jzLQFkvkWP/IgImWOuQj55FlvXEnmo0YlHa2snOTMd73K3bri1ju6wZvzIIgtPXhu7qSJgMG
lcOVWMC/754Fpt3HrLYtB4vG8OMdjdTsFQvmk0QIg5RydyfuW9gGW+arlHFnE37xqAKeSg9bSPsd
S1BBttcBYl73pAgcTgUtE24iAgiSs/3EuTOrVHgiW6xetCOm+WRJ59zH6pO37hFPAbvf0ShAFA4D
L9/nDe5z5QswtkCLYUcYjJsAJu5z2/ytWQTh7GaVVIhjsGwSiJ0A/sIZ1sgHOeaZ//rW0PZQBVfU
RB1ZDFyc+dA0hqCXM6DtK5fb6f9ML/Gdak3DtArHseKjB+73fa7xG7LrPH53E9yQ94XMrpW82oCQ
uZSRLbC7aw4AimbcLtGRwe0grpGZV7/2xKiClFrorkJzFhs2EuQZon0zGaHLsVp4JzY7deXC7Lra
ZSFDEcU8BIhf7lv/5HyQvHzyY9DncrsrAeA8Hdx6Y8/bpiemIeQQSFP7A8NocAODv5Un1ZyWfUM0
zNp7+BNjqIooLhIh5Q07JwMWegEgvhAnGjqYA0wpNEGZsRqTJnRjmlDcUcfsVNWsir8/RBxhQR5c
RjNQ7+reojE0PZXKNt7xX+e0gu9gmZwB3zntUTcMGFfa7HHb0j7qNo4lLnrXEkAZ8devrN3aFGDq
7L48sIST2I4rrwsoomRdh+MxFMt5XteTp9na2wtdTBXbepjRx3YvlBz2mj9E6W677HzegKXXxzdR
uLrK1rP7tV2gMju4WYj88tvDZ1gMw0nzctXlAZjcuPHr9np7J+ucrXkGrHc1xKaJVYcSzQ4RPSv/
a+aTgPOS/hWgRHg3Ez+nH4Cjts3Vd4ln5d2FFVaobfMzpqZ4xqbwxsab678GPxzmRyTwCN2/675U
MTCHYfurs7AC9fvaA3JPxhe1rVHeu0NBZ6kpWG03JosfHWs/iKKKvAeIMg11BQVZnpGsMfVuTjLs
GkLMI6Durs7cxGs1RcVOSRUiLkEROKqV9xa8+P2yecnPnK5HhwmKWEeAcEQAyexNnxxjw7rYg7Nm
UbX+clwoExHHryqkv6tkX+aPwygrbGiFrI4vnmLyHtiJaaTGPAtaGEAytx5kdabvt8JfuPKew3Mk
FB9txY1xTbIcE91rQtRF1NONCLwkv0mSnesMDAPUqrLlLcKICuuEVokE2T7/9BlYgodJvx1d9t+d
mqoh7/MuXSFOkHqV5UDKV3BD4hKUzgJUB+QWLYZdZDaLrRR3LmWo1PPTU+hH/LIi6pOvjDtd7RVW
CYwG1KFhSpFgPCyu7/wlcmDUa1SznbdYnqF8VVJVPZWj/knNJfybwnnz2IwKvmJBwmsXqSdBpM3R
jWSGM8dSIc5d9Z+ra9qpki6+0Rjr85N1Kea8+uJiR2IbJ2hXDjeWBg4n8q+ymjyRhvog5LLGIuWl
/N/+lzazE5D4n2aC5G4KJiYVXxWUOaVzx2zLoihSd+Gnp45qiL13XBio1EYpIN0b3YwPdKcT7Bj6
14OchcQ0N0MRXr04IfP0Cp91OATwAVu1rWmSyEtvN0s2DeOY3ZXNXTHgUF1AjrniQPhD5rE01/NF
ZBiPCO8EhjSnSlas8+E8zBjUUnskEjOG98e439xu7JwX/eJVz+OGFxugDDoEeqY/MiZKHk3dRnVM
QOv2KIZaav4SEvlC/pZLBiKfGooLm6PcS/cORr93hBnzoP4lQVK6jz4iu1WsyJqdRStC0WmuGJHJ
w6KxYz8hQGrFE/R+3ON5XWtSduYDKQFipZ1aPeqNleo3HUloLnEKSggDS6mUEauxcKNzcUceghsd
kPyvjx5XZQkxv2gteZngQwKPXDcPHfgE2wzEEUHEbiec1UvC/dRCSlUCt5PnmLpagmijxDMQKhOK
Kmj8JxacvuEIpQlQVi5Chmu8fBiCHB8eHUNCV/89Aa+BSK7E9xWRJIUgrYFN2wyW2JggAs6fLyO9
pQNJahM9HxdQLWIllm3qlq3rwWZ5caSZaYfP50vkK/7okc4GM1tOCQ8Jnk+QeudQgVeWdw9/5rMi
blE0y5cXgPMQy3hfwcfJzwsG0fi6JjVvUf6an9QTf4XaHlq+9Yj1qh1O6r8wcCArbUsT/fv2dOLx
HGrSX7rA2bX2VzE2lA0VO2ABkL8swmLY1pArz4gfH4M25fOjPE1n2T9bDEooNApjL6pfwlMTPHXZ
qJcFIwQndkVRQbwjvFuMv61PolPRflgPllGRqY2f9iUza1DyBE7O7wCkwMypPNfPL0NPiytX94Qh
cJ9pnSU/LeOpv4UT+ZK2PofDHQEaSwwenjG6RvNFb/hgiAuOBDw87JOpZadKeF2nBUvja51LfM+p
hRxQbwK5cgl2nRdL9PRoIUKjUfKzcKz0dwvZdStiiCKFlmXH7zLCd+ohS+3DE3e9njoGeTIYhoTC
MObRmsIE4IaRbOlR5K0cDnpi8e9kda4lVW0tao0I9BtFKvJS6Rg7f55JYKU/sMFhGL82ECesUfpe
grdDkZjtsTx9dX0Ha6rgENB/v4NNr0V1J3PaKrEpJR/9EhAjP0KVPPHXy9x0Bu8vLkwVqk42wJXH
uvWW0BMtbXWh/WoQJvq/bfwsU3S4P+xffrvEU8QtgEcoPUjCSKrE7tkcH6IY5XZUk/sA0H+g9HxR
shuh7e6vnVyr2VT0jDryHQunO7Xx5hGXf1bSi+dx3MfvUuZKewGutZPdmkwaX9LoYult9hAIMTqB
kqWPFHh+E2UQtA2XZ8wVt4QlqOLBQGttsNGiizKVa6p9GDx9JZr3EDscbYM+lNCDAKOJtmaIKhMW
rvH01eBbNgd/HU4RPqNftIXPsQwrz6Fyvvq1j/V87hu/PWjRC+GeCDIba/gsjfrtdY0XAPe3lSRr
ZtRt3FH8pGtF0b6IMeCf85ZntbPwZymObSABJgI04drIlDb73QAnpAHfHqP3n+f54/R6nBCHA0rH
CmCsXex0lH3km277mgt908o+rxdJAKEPBN0mScd0C0KG7228caeaMUg9SJcpdAWKyIn+rb+0UpYU
IcSGYCFM44zPZMa34ySe/Rn7cIeq64qAUQZI+cD1uZdntcd/R3oEIPSUlzdrMF2rPNHDeTL4Dbdc
3+iOSnlop0W6YFN0NxRVZlYU41/yI4swNdSp2McpWcWhTDI8d1bPxTjMjLCk3Y3xhvZtqd1NnEYk
sINolLwfAkwdyUEVVRfoPOQKoribRGbYjRQzidJlbvWiADVuwNqEW0LNNH4BEO+19L9qnOxRG0eV
6tJykkQqx0NzI8kafr9wuTSblynAXDUu89LYBpT6qQCuAbKSg3o00V1qhPWp2o4xS15RoYf1R7YL
52eY9ZBPDqhVkAYZPJHH1TWnCK0ekhwhv7lEty7BAIG8cM1+IlzGXZkTfdHsNjmK4L7vPG9l2jp0
htYp08O4PHUmyU0OeB1pi6Ewu+bH7cQ4RTZ/i/F9RQSWWglYk+GWWAYs7/fKtEKpDFdAj4xar3QW
kgxHMji2THz4VVz6u6NEtvNxqOezSy6ymBhrBaMIwteruXtW3BRqMB7DLYkVW6TMNByCbloIm7QR
noaD7qM62a2nAJQ46HBsYtZ4vdOVaYrMkE2Y7L0nUogbt7lZcSxK8X+XKnfAl3liRLGZUHIL4LNA
LIw8TmLxN6Sc3QG8ykCfKjAuvHx1x+BbVYH114UhZ74kzUC+E3NVLtlmmiL57JqM4r5DLAhYG154
ivo6l3eEKgYFJTYbWBGjCsD0yr86hqag3FtwW0ZCpVHr3/Mp1QJg90sTNsQgB6G+VV15mizoQDWY
SqxQVXe3+G6cp7JhivWfWpGuSIDswQRTNztQRaJ3FKkP7SgP4U9d9OxEFoxw+lwXudGsvxR77UQv
oJZYXIn2YlNy/W2+T+dw3mE0qwTaN3RadBzKYsbmLNG7U9KPcXXM19crpepbCcDGTbJash38/Tri
wpxuIRjIOvvwQUishV/InTf+KYCaZ3ZueRaUcwWkrYaZjsJN8vMe+O+LP9vCNWd4VH+T3U7sqDIz
w1t/7N/S+3OQJmp0vvN3IlxQTRhVaOd5gmbBT0RZpBwB4LtBejPXyT7ymVVGEV+oB2tvHR0VES7E
5Ba3lkqU7OJtie7fG2L/p/goAdhKs1J3XCv+mnDG7w/wIKRgoZ+ewUUqW4wHhb+IiW98/uzSwEm4
j0Kc+C5DwlJrgQlm6XwuOkfLPwW/ysFRJt/rHatoMLX7bUGj42iiwrQ2SSnDQyLVlbsQ6sOd//GO
XQUyqt6UDAW5Vf9SGwAvdae9700Swrnxq3l7WC1URuFxWG5JkF7cNb7El/GpKwrs0xGW6e1JM+FH
Hndzrb9LLEPdgb8fqeq7gp6m1XcZdhQxhCEW97kWCE2RIPXw5RdCkVA5g0ywSCPLWW+hdWewMwQR
0ZMNTcBNiQ/NE83VdmJRNSh5OL0xY6wAJ92+BbZSMC7cAvdYukKOz0tKzZ/JhSWWF/RfGDrJw9N9
5rlfz0aT36y19CKpHqpqwf+EaXQIOd2lTuDbUivZQ4Qccg6grVNsO/7uSmPWk6JFmdOVS2EmX4xl
sZ0vgc9IfwI4efAR00mQXOEJwdaU39Nu6aWXupxavprqJjiAtxIWKW+/dfAFpjd5Sd0dA2O2n+Eq
EkLVwC4slAmMDwKNQvjTRJZehdmjvwUJYX4t+Ac7YUXfpDOwabjcQpDdUAik0rcyV7ElZGD+5Y++
EDwnMegA8N++WzIoIf4M9+0xoFGsqw9GA2aEyrdTUXa+byj3JbeWp7ol9lxwPfBhZ9bG02ojFQia
4VzklyYtjTE8CCfdnfm4BARQT2cLMVwVH4vSm0fWIuATXyl+4PnPd/CT9+mNM3BQjZ2agyyIDkHX
x5sANl9XdG7gW6naic1eIGvCqI3ipkattTuQjmeCMauJJ5AuVp4rzijDbFzfDYj4qAdLfSXpBffs
V3vA6aRRUBpIBVZO0jKL9qF9R7xXiCkc6L99zlUApZECGaFCKK7HOh6i5xYHhmAZS6R8wlDhWvg8
0nLEx/KJ86gLhl0A/dhVX5jZzsYJtcQcbshWJAShI3j6Swxlxc5QKNpTMf8cSkthuJMff+YBJIpo
jfIz7dR48ytZR3JRZu/wWXfYP97PjQt3bfsoKvy+oSBv69JtXHhr4ZMkR5xWtJXCqIIUIy3MpgY7
M4CTeqx5GuFD3wFS+/3KCg83bXO5OUNs3aZaUFOT5/WPgPznIAmygOA6+N91UqmS68FtDHtS2uWH
GVCuNyKO8TQJUMVFCFxs/jaCXwHKe8enbKYOkUXBHhhODfOsGnQCtbDnLx7OxeZGRGLqJijMKzq2
z076tExDlmOvojUpFNDi8e+J7uKL7ym8WoYvIdKMi4Xm7qydLmHyLRa87eaH3DG37BuXnnnWdz4f
gAkZ1B5o84j8CJT7LNbSnoBZHmXlRcT7zvte5KlltAXZwYLj8vh9dJEKPgnpwPEdD3dC71IKGqwz
H6Fg5ncrtxl/o6ZXdlHbZuDGzCgxFDObnPNrka1Ws1kO5HKrG+wBSsobbNKS5Qvr6n9MUa23R0ag
SsEJcoM6Qo1ZfthSQH9Xk/HM6NrxFj65bYZCkvWTUDJ8RygSWSKxHsFqrIJybJAltWrh8uMJwc0j
ZzfoPrsHD8bvcBD+s0rOQCYYJKRmv5MNamoJQ4xQWgYzWdcs6MPZmohEASGrwV647sW2bEVUV0zB
NxyJqzaZqqK7MfPM4RDWDKMQnc0rqu7ZNRPPGAUw47wgUxgVSXs7zGj6fgze4KAs67NeAcVNR8yO
srehz9zAVU+5OBvOsxme8Rg6//7mROzdKcTQL+4uYsvV/i8FTye8ddX/ayTCs3RiuGPU+ft2pEF+
o7srSVWyvOm6o4NmIERb61KUsd71gpP5JgG3DSgusKm66jpOG1IauXh8fac6nt7QEp1Hb14U5fXq
Hw9oJKmSJtMvPR+EbX7kNsyw3dHyk7yTubS0dVejjYgC8mSGW0OAexvEfYOgipc8XcpkK4ln2cuv
8rq4dtcdC0orZ2clnFoNtrSvuwTziTVCgGht0fK/98H+HTrdH+Ttcv54yMX534lhfyNYkFxSLyyO
knvqRsqQLHViecngbEQ+0gXrxb/45qT45lVVgiKzOWsW5Oa8wxG/JP05eKk8CSw+cVSHNTgatI6j
E7X4SrmX0vy1aIKipmKaZ4WK7ewRWBpu6g+3WxKlNZSbdAW+xEbqUyXyLThYv9/FQkDqJK3XSOMU
tAtXEriPrRxLtKG8626Wa/y3quty0pugV62CGHzypZMeuS/8czuhkV9VVixVeH9vx7MtEIKniuPH
jufu+AOD36o+1o3YNKZ/4/80SL2Hw7kW4cIl8emoqMzKb8msh2qEQhYO30+TkHIN3BjlE/i4RbXa
Y3ayRHk0yTaayF2M+yTz9eD4ajuHQ8I/O6iyuQiKAoRurmO0AI4duLw5Z97ttKUnsDR82Tu6J4k5
nUdnt+xodXS+i3WmVhOMu8PpnLT5NeWqSBk34bvToWL1P9Mqa9HlrK7zf7eqRxnhGZ2CCopK2ayT
pESDW78mHTm4c4oaQJGtjZ2DTfzw34eoEVZCYWxuTgadGR3FKyVJ5nH/FjlWzVYinMl5MvV33aA5
h7GBiQk4g5j3cW/JY4tpQZiDt7pLWK1H77jckZ9JytMelCDVkO07OY41i8bbu9q2nzYznfmLjDXu
U1q53xWnx3FnXqv+usVoyZRqJ8Md07mDTkZ2WNhqXd4GiROHUoVXcr3u+nkmi2NJbdyc5GAZghb4
dQDoDYy4dVF1Y58tZCIrXvWeut5Ms4VeTY3jqzqTgtA6sQZ4WiUovbPZSWlndJo2sL82NpWr4Sek
4+cxyybiwbTZ0OYa/JIR9usyYxl08U3gK6xlO7U5oY8GaBzy18MWfqMUPtCvElvPNZKSi+N8qqhj
nzUF5vD+voIZ77AuVZ1Pazp139dqv7+znDD3mQM03wUqCe/YZOvcexHz+brFDM5y+qn9b9AnwwYB
AWGIfP+SsuqleLVNzbae4j3peOIjgnDesEbm5SbAAuyRT2ktGkaiau1ABunpga2kxmnjLHOSARnt
RyxitaJsrFNz2q/9Qq/jWtH9red3Qx1xKcinQUsjra1r5RwzNLM0/zVs5c9+1haXhYut+JPJZePd
RU5TuR+ZbLsICLZw9wvb7aiAfJLEnljAnvoCu+TwccF9NzllZvD2EYWpR2psTM5c+IJz9S9KVusG
qyt+fwT5cFQlhy8ofB61OrVtWwR3FrJhDSfcckOhB3Q7MRzydRNsQhyRxJ9TkSpZQrvdu8SvATgf
v4yWl5Mxjv+4AOivRGpvNFOykWfPN73Bv9Gx1VcZgaOdu+8m9XvPL/lJd9faEj0HjP/atFEuZA+e
21BE2N9kpUhQCs4XI9CnEUiGzF2a+ExQW7CBQtBHwgcwk2f856W/CHh7yv2GbmuYYuUci2i8xaQ/
YPn2ZCT2IpZ+JgNxgnMt8Tulk9dEKsjmWpDVNo6IILDzjp/JsUgQDG9r9fbouloOFrdZlxwSC8Cb
bwm1s9DQ9sMn+JYDYvGAv9lW4Uy835jaDrEyQ+8qNo9ELNKfIPQ8RXYbStt209ADmOeONxjsIfQg
SxOFhrZqf6ldIfegHdGSUudw7IkYXbEVACmCYUdqmG8OT3EHC8p7ECONvzYgamgjpsnOWyLuflnw
K+8A/lTuomBV8NEeqkBIrlT7lhaxQxm7RUqwl1Pk0KGMpcW5cYPirj5gp+zNl/YRw2rfJl8owB1G
gqRwdw6zTzxBgiTE5Vj15fyExwQ6pQnqPY5d4RrQVx444n/NijyGQ5mvoPh92jO/tUWQau5PXvvf
Z6axWvje2FVyAktveK+3cnGUmQanKZBDjT234TM/axG+43VUD5eXOGV12og42PQeo+NSA+bC67vw
AX8RrsBLrCklLRkUqnW+Rh98cUHY90bH5efCeYdcfcgtEn6rO95TKVLlX4CM6vx7rSIgwmdzkzYu
eVBKOGOpeUFsc9L7A17pzZP0a75Ah8n9JGF46peYlnHboxO2qBCwoFVUU6GbXRvTKYSUFc9dAm2Q
T/fCXofQ16rJdNQwZSK9+zgSsroh0F6YVXC6h/XKMUpamfgThN3waDhHhbIFtc6S+Z4RNHxaE6bl
Mc6m8W4aM4bTXGC1WGw9tdiC942B7UBs7AmM6ULgNogXmhZiIkREmBi98q77F4DKFv3CHQg2/CWP
HSppXCtIlaZ48royb7PgEyqby3jj+QRyaAkWyLvd/9Nzc44lnzkcnmZiGANDmHfm1LDuC42MRNUh
d2k9h4KqpWwCRDR/PWzqjwjsv6shpz6djyiGEXGug1uzjncL6ycwcBZzFEwGhiNQTnzyrRs8QqjS
hKfe3ssbiTbwVzyJM0hae8A1fowqJcMY/tkm2swz3e+f0mzH4eM3XBNaWJx3NfwJ28Id0qAU4S7m
EmKFEW499qzJNVc8Kv1dk0AunfcAUrmzTEdHqhXuqz6pOYAg9a8Hf8YQjSn+OCukz+rYdtxqEaHB
Ha42r6xV9sUfmNNL6CstuNpt6Qfa9qZITHp35a2bSLViyDA/es3uOQwZzp3o/ytV18K+ril+lp5R
EVInb1eYWHQMh+QKZofC16Of8yD9bYtSTUhpDxbpHC/+zHaHJSU8TeYEwLjBN+OgKvnZAucuJvBA
JjWYK4vv1YD6qgz7Lmky/xmOidybN+oaZW/BJQzfALMJBzBghWv8IRyvt47TxOZkaAOgRY+e+xnt
qGNxQSX9wjRmZFB4dcABZg2/seLNBRiDNM+JRTfqxdMWYiCjw5g7WMw5zTvo8MzdHVUFXg4fCLj6
x8WGFOoDcUXdYjrZYqGevKl+ZZLDmdhb7F25i7Sq33cvXWVVEVPPGx6jMvN2PiStjB12t3pfOvxx
BftFlLyOUM87Tpi0szLUR96zZxP6FaA+9OhoJo6g2WzS87ChxIcNc0JTUmzltVTECfpIy6RMcVHd
1a8JU21gthc3Fr60Nmozt33uKaJMkf27bk9GlPr23mtSBQo3hC2J+gxIzCwM+u15udV0sjCrHeCQ
YOHYHHrrKpmUjOV2r6mIpRpbpoHEFU6s4+uv+19L3XIqErlZLPfsyq/Y8wCnvebyuPjzcvnegooD
SDqv8Hy0xpA3ryXJODsX1DVnELMB2g1mibWhdn4+svVs/HZxSQyOvmIkMgeIuO5dopStu9coGZed
hhl81J8jR/4ffR8+7gKOV5bvc6A5xM4ei5AmR1Rz8pBllGQPECVwZBR7HQ+Ihca7TUHR9IehlH5y
FQD0tX2Q8ela0gllzyr/TV0omNUE0uHA0UjOXDFAw0GRSC2oqtcMmR4Xz0aNkzlq2q4uIJGyXMvY
39t1xs05mJbGO489/LS4xL1Gm/7pLcYJfqKD1FHl8m8y5KIz9iFIhS9TRenqOwaI30eOTtmUMJRw
4cvVuvXMuFbb9Xt24qTVodwqPVyy/1ocFpiICBanPcypXfoqCpZMiJ3NoVsTS/+/QPUnTvJgg4I7
AM3xlqJ0AD5gJx1sZe7rFCRj38Ui4Nh6CyI9l31uvYIEhdkXRD2ILmNaVWyKTyITAB/l856afdlP
zaGLtjQKSwq7Y/rswTSiSn6tN/kaQygAvQCT4OcxmnOcSyrXcQZncNT4VmNBEXdbcKZGoMZXZgMq
xl+l7E7IjG/MG8NgMnxE1ZJTYlmOu85u+tmCkPNR3VAYvGR4eXCZ9Ck4BqO14gDZuZ6XqpLTeyQf
gx9IWgUunu2ox6j8P+ecYuRyzap1xGObsR9E9o1jgoKAYhMIC7xbzNuAY9MklLzIVVk0jrRbTuwS
wigLmnwaNI9owtx5U1CGdXrObF+SlNcJqFY+M76b1JzRu1HGlj2fVA+bYY6nFSmTU0kSn4Rp+HlK
dCaZKe9lom578W8YKVaPt68YPaMFxTYfaRshjBphDR/WiyJlE9ME/JD0D57EViPib3avGLZ+gi9D
pJF65DdVO8EAc3zH3XMBg43jerxbg0bFqdHLbcME4td6yaauOGYyn6BqsA8iKOce98hlXWSYyXyA
EoDCGkvg6ZXZ/OmghmrGtg5swjs7849No9OmfTDgzWRHopQ3MPZ2oe+d2OHlw9RwsYEpVZ6k2P/m
Nc8Kly2i0RLtGnFNbR7ZI18Hgz8fOh4fLsVvb/Tdot6y6uCaDG+3ch+XUgmauLgXNtYfHvntYpcM
lzp5+4+hV2gyZs4Cgy21/Ve4PpOEW8zD7gOspAp6QQDO9XlKWmu4eaTI9EiFfurjEufD3XG3DYo8
lOrcM+mDPfKnpJ1Th1AlNPiyJEAqQJyIYtTmwEWFwm4+tQwq0NojaXyu29om9yI14S6bHx4nMhrJ
/ta691c0IdsTubKxz1uKIHmAwAWdf2gf4RLCxr11nxflrEmCxMzsOA/IUW9usFNZ1ZSYnZibDsHp
u5yel55hWR03Y4IcbATE81tEl3kLH8hNCt0xnljSHfZ3mKGH1hyVSNk08SvMwmTf0kRuWOVNDHe0
NmvwKCrIXwB/bXehr/0bA19SvhCAPsMgvyZxFzILc2wjNqaQGphMr5btqCiolvjpLNHIjp4S64Ob
Ea8sNd0zEd2WFIlxY578Qc1m9OjgUsAorymSpucpy04DS5iZy5F8bKaWQHinvcsPAcHGyCqc38Yh
4mm0XvKDmj+B+OQTFpZ2DplDezRAEe1pu5jtfDCa0xpQcq5w68V79u0Ca3Pqxs7VX06ej7R4T1xR
C2bctH8+8rgu1HeIK1jS87osTSwHOcu25aqf3ce56piw+9O4kyLUiWb/bXQiONVSOyHK6CtZdpVc
E/457tS7ovP5kuS61AOli9DsKJ7yTBQ0ro57/28lx0HT0q6BZgNvBVQDemIwqvtoAV6gAz9JmXN4
D/Y3/buvLs3LsyIpImftb7Y8UB6HSKlXwWDJuYz7bRxPJkyGgxJ1apb6acB1HkbeL0FLXfRkLbYc
eJNE6FBl+7UDGx9ulQzzOPq3cnHlmxSoQ/V0fca+9ZsLwDo3gJtNjJpEJpxuI119Vo8ksFlwj3U6
qYCWWbilvmg0KOVi4kii5/NbmXnFZ7ehz7mKLdccwUdQ9VpnpArqI3r0qoK8rVl63cFtrVvDVVyp
Gm3JqNjXXtrGPDNRxBkJwIaFg/+42n1xSHaEmRpoGJb6norX1nDiKwkc15XGs8xUvhcmCgtlGmLX
fb/5ltEHZMNM6l+2ApVY4GgZpNqkG7nRxnE6LL5Kn8PlGbWLTpB3px3Ekuo6MLKh4zqJcPBgraS+
twWkVJES77M5SJXdEmoPzZlOhWnS0woekbCJndKu3W6siQpT6LQCSxaQ0NUveqaBRhyh7dGSi3j9
N871fXj7kI0fvsDSTEJDoyF1sUT8dzCBPgiXPuK3igaEIfpbXue5Uxww+Slux6bmMpb9ZSeBOYql
Qhl++mOMvagR/aqW6G+vpLdcfvD2Hw+qA+WnySdilnJuFX0N95IKKX9XngBvCESFFlzqxwIMb2w5
GoDclFYbqA9E7gKX4jr/+NK5q1TnGkjE+wbNGPvGHmTFcINd8RGDQhahFoZLVhfXx6OadYWHT3YI
fGH3ZncGuBoj0qV6DmTarS7ChwhhpeHJyydFSpJY8X9AMB5bA5rPo3Ti+s7RceAKfmxg6xthzMuv
XJnlTFNtWb+eWdEpa4dXa6JhQeYUcrrPf0upTVefmTJGcxANk9yUe0O01wJCBsAuVedbIo0omNqW
1w23lTpNaqyVB7jV3RQsg1tC2cyn19sb3mF0wXCWaMsXpkNvoZcapkLzlXzBWyrmSaZRiKyTmU5e
0qAtFFpNDiOLikMJ9GTfQOvC3kwBTSSS/Ij+WdiOiUlevJiZEphUq27OpMTmdZeOIOefsEE0d4VD
ZGvC2cdk9ZGta4LzziAylGSZzT03Ejt1od1MJdjVlc5lVfeGPhgm2xTUa9OvhivziCu6Pl/dt9bd
tIl4YiErsSjgiSJpqBeA/Kl+gVnk8O+lp1cwV4IGzZb0me3GpEWy8C/cgICMuXwKTsZLTyaNbVl2
P6+WDJ6UUoI562FSH8PTF0Mo6B71QGDyCqptpZaL8UwyhBtHLOQkhPbfbkFkuzZzgNy9cZeVy+jw
9MRdrre+NiCDKQv2gsJ4EQQQuVlvjExd4KSalJsUdTjKe8fq92kmtz4BOC9N2tG0sQwvmQOExwqz
wRKi0F+whCGam0aSosMMgJryH/pUOtf8hIQfGYWpR+GY+pYuN/8KzTyFeiHJ6EnJuk0d7Hez7cjG
IyeAbu4TrsZb3PVvkeAgkBn8vT/2NUqFtN+V7voly9/Hl6d4USQ6gHq3IRxBHFXAjDFHdWFuEn5a
K9OsIeNV+q4/Nn2VjoC7Jfqfx/lXfs8cGe1EwPXlwVK6/xqiL2MhZZ0YvQY8j+BEvhFf1GIDmBSW
ozGMmL39R5Ym6K09a/13CKdVu4tAM64dX3SKi2+n8837YlArbkwjtzwhS06OXW5OUDLbDKUzLWrU
LzuY+kLI2iA4XM+B4/kv5ZbZUn8ecYvBPjPLDpfur4/zEGg4RciD38G2hhKEY7L3QcIuE0xKFrTD
ff6qVeOiXx//KE4QuFN8OvERcP91aC4At8+Otp6rWuNhAwLszMRhW8E4dNmC1DJA5pkFIm+xlC/c
HXtJ0UjwombIVc0gNRPED4EEuZ2wa4K5ontq7ueUahp7r/T8cgAgiG3iBrb8W5PhG1JpGmcusPqV
/X2dG01NV6BFkGP+YbiYUz0vmxjASN9feDRGT+25VkEPLdiRZsaItyT64uZZv4CkumUQmHEd3t5V
2AL4l7zqyveqnftTf8NI37rhI1pXOLRpX9ajeWuxZkB7TeBXS+DrJWW8Shuv5VgO9pitIfgi0Wqc
Log7xuOWS73yB0/wu/tTZEh2fr+mR9ckpkSGQwvsDVKbx4iovJ+F0F+ct/yh3HL1xu4Qoa0Zw3hR
15lG6QGuLj06ogtl0GFXngAHJoDqK9REch4rVjuYhY3glclXZ4Kr5Xvc9mUdqhGaxAQQBBqRc4HZ
6yAAUlge0t6Lyc3bmL2G/K3sN0qVUuxJHfgDEQ5kibGbBZnGAjTafXcbVJqW7O4HW4fAdy4W7lJ/
NiGjwz0zaSD0Lz0by9PtiabaY46V+38kYEN7V2+YKkL1agTuaYfXyhiZrfpWqle+9hZGtbFnz99v
I66VxMgcnTIUO2GVX8bLuVekI0e1CxS2U6PiOBBD0WXVrQTUmO72onH1rmpIXAtAUQiX7iIG5JxS
X7BFmXiun6pTcqx4AnFgGgLwrXf+17LaJsBRvfGHVrNk5/L2OlJe4nPfHWyjSYTwP4q/dMnz7Oaj
71ogvf5pe2vR3P76GKMVJv9tpMBLVBDMIy8wg+cDkMC4NrSH/notJqKhFm5ObEcuWSJLEX8yiobP
wWZzVO2ZY9yhruWxXjumId5gbp5xhqxVQjC4hk93X9giE7Wrl7E7q5IkgdhBFZ4Brtcv4CTHGeJH
bYUgxOoskt193dn1wbB+lgH/3U+tX2tavham0QXz187cicFGiemMAY8owXLeGcpBb0+jZDcx5hVM
oNI67BsfTXKxXwB1fCG5GVKRvq3CEyzDzl5buYwQzkME8ZsaF0DO9B/QjbaeDVxp3ldfNO62slz0
QdU1oUFHmrFOZvZEZsgkeVQZHv2F+ALiYWB1EPWKx8d+mU+Tc5p+pFL8YCyRHEjK4YHFgsbF/qhS
tYlxh2lICyykimipOC0cjcN2Nck3bzH8ygn5XI8wGZP9axpq/at7E4gF2y9oaTG5XIJUT7tBCj7j
G4lOb16aCESDbowAVOUBfWqOzDejQohryFTIGdxMi5EMvBfMqOJmdwc89D7OsU+Wm5C5mi8171zj
uz4Uu64lfWOvNyJCOaE5yRi+85QaAglCI2PQsltYd59gcn3NWHjOR/vhAVfzCIxZghQWZdbmmc5o
sXiPIy2govB0EC1/dFyLo/6xOdPxry9Dfi55dDV+LmRXkiN5Sv60dysJn0q2y89ufJ3EFjp+wzk/
DpGgq7DsEPJV+ZrjLM3aRSZxA39tRqsaixvoyekiPPndyN2S6NR+UYdpzIdoGSoQISACNfrPhWZT
VN5ocLNkRjc2aU4ZuaABbSlPJScUn7/TknsTD+3GjkbCuaKGlDt5YfoV+/cdk+5VHmW4iV5pEG7j
3oB7klMMHmrHZ324QEuIHk4DBlQLdXBfxzWGUXcWQp7pxAPr0W9SBX2oD93oh7PmR8Km8m9CcYcn
EIPuB+84MR3ov+WB6CQ4h+6FnnNcZ1TG/4sUGiAwhDlOKXhfyyaCHAKxr2HVbm8N1aUvRZuY0RUP
pBqSEf4qw6jFJKZS+KSRL9i5KpoUdmz/kMCSqPS4mgL56Gue+6t1KQtNUUYH3ViHf1RawAE7zqXO
z0yTGafIbauD6ByZq+TKmbhv00fgj/EhJJP4gNMO4OKaJxloKi0V7fVyz9QzLnB/uQZvyvdpkc6t
up0/eVEYx9Z5iD6px2oDtZl5UGs2xYyQ2kT2lgdxY1+G0QNN6m2nsdz1BNUdH+ZasSgq5fTZfnTk
/B8qhwDVw9flz6PCOUlgBUVU6LrbzH3+GgCItooBCSlZyIbGQHxO3ReR5/YUsJGNSODZDbbmIxGW
y9Wj4/dOglHTqYju30qebhTmFsRDkImn/saLUMHNb+N7XgOnhGWTg6LzpLdt6OJcY3RviD+AtW3P
5+wDayk0ilhnksYUBs4XWAtz9Goxm/4JVzKUXl4jtRc7nTgt3TRolGYkvQXr7bdnKZLa+uKjyQSP
E9ug15tQidqfqfUZFTjuxRo6Qs/YEa/j6Y3GHNlSUQ1I+HCUfxqcLpPo8coutGiQx/J9G/o6EGdc
aGa5R4hQSlh8X1x6limckVhJA6/GPdsP+JovAxntVpyOz5AJ5pUbEcLMvwSEXXsoM3/Z3Gsl13cs
3OCG2xCTjukuriafhnwwn+MIpQ/kMPCWoK2r0/W4f6UPIRGjRxIbAwRNhQ4R3ZiZapskJjAprPuz
K7R/VIqaZNMnGZu0tpf0dDgYmCEbKufKPkpypim9yjUUVxMXPBNIA5R8hq7yHn1Yjkqcra5AY5qa
YtSkmmR6UwV7bogvbk65l7CMcjQ+q1REKI1NmM0gRkqm/T1kNqTQ+2XfodsKbnReuQhNdA7R+5gA
F4ZlyN4gnVYQLv2cV2+6s+inS8/vw01IIIrKqQDmEtHcKJjgjXKIYsdzz2481f4eiT2dzY0LCir6
GxtlYfCbbYuDg4ys9Cstd73Fm4YzZvv+oRfiPcJP1la0D3KL/N0O0qdGvQC/Mk7YQLN8EaLTXhZO
q+dEWuzp5/pNzGeilE/tJEEDje1Yu0gN737ayJyN3CcJH+G6aLOoovVWm89tni+OAs5EwSQmFB7w
gFs2AWe/uJUAt8F5TCA2uy5qX8WscmoIKevR8tYVa6VVqofhpLEozyCO6d+Tn/JUkN0Yf85+vEcz
PQ9lsjOqC3BFrkx3carpm5iz4Wc2bp9MYe/T8S5fGP/vR30DzkzGnQXsjPuBVPN5qcT29AqE0I5l
rK+uJuCmvDKRaVlTDBkyVkz7GX4FxHJN7MN/bchvDlS3WT1LpgWA6/fBjnSr0uNIS54cFO4e9zcN
pszAB+vJWilgie1i5SScG8J/HOdtD2XkDNCLiXrD9tM8jEWfAvpBFbQmwLHew8c2ywFtgHG+6bDc
6P0o8FUEY/3aVGJ/cIc2+xhrUD7izhDRQ03BLpRxkCx1tuN03L1cB0xWMl0QPyHv1qUlP1qYOsw3
ZPE9N0UFzUf1Z7Sx71nGQ0Dlt9q/9mxH9PTAVIjg/ljc3p8r8+BpXKMSEB4x/NQSDP19Dk1Jf50i
drNCicbZqnCZ+T3TmVtr3HUPL9z/HrolcD6JxE1vkjZ1n7D5czXZ49NlbA6RJlIPSA8jHjHLMj0a
gtQJA9ucrY2forRlNT4jly/hNdWsavXC5P22+PceU1wPpqbaPYx4VuJKTstdFld+bHUOhaiUl5cY
ojurihX8q7HhwZuAGde7nC+YqjhjR+A1H6NWN8jBeMgLdCZxqOAHPS/hRPgqO73ntWB7RSuf6LvR
sQavjyRGlcHKKKqeY++Pzp+LOleKtgwHAZESQ1zNceTFIEMiL8xKz/4UkudGv6pRJVe2BhHZRnlg
QK0mqcZ0hruSQ9At2R5KOt4QPP81OtJT1CMUKxLsATlyA9wF4tI3hk97lRxoTt/RVOHHJsY9MSIS
V4JvBeWbwWgAPjArInyksS9hNbKOiiVZ0xOv5Nrn8f6vc8RsNm9r63dpV+H7VGeEjA9bepXeVVg7
Z9lwZRyDAeG9YubD6BAqJgExK+jLYRvfvPJC8wOo5/fblUNCEx6ZzZ/z/c3uk00W1imIMlTuRh2M
W0V8JTjrW+YzMzG/RuTJ5OO0EmGwcnOnAfhORaplJG5VI2Vm80rTYjrx1sCze6iP9rSVEfriepv0
PSf68UK3Ace4L2X2J2CpJbJvZn0fZo2XwgCaPcwiXgg5DfrA4pC3LB+VNsrCDpO8tisDse8d6LgO
VmbR+nZJ6mlgOkatJZfD63ugyRyffbn6np+jesGX+llh3LObGpDwRjnkJg3l01sKlADBTs5yMYsc
tzWf1U1LtablW5uPyOI94DFg626JvDQEOo5B5HJdajrEQE+341AEZEgGYE1deFlcYXR90UJFWYe1
V351vhKNZ8D3HQORVh3vi/xzJ4oD6oijWkS5GG0HRdTu1GarUccJ3G1S+lJa0a+9ixDxawgo2CZe
M6rAFe1Bmkg3Ootc1V2kKxzKL8v/5Y1x8DqeSy0WAPFTDB3RXi9MZtyDuqub5GHlOWVZ+O8HvIZp
aBlyCAblc7C4R4ipxjKW3Xxx2qbMooDBKBm/Xo/cTzOrmKOTAhNPgwaMnNqGr11YdhYE5mCneaUF
k4aRMwp3O+Tqx4Qp4KR2Ipc7qFHh9Hw/C/SUma74GEjYvsuqhY9inQcAIB31GEQw7DHe92rwztFI
RmUrmaHYednHq0u3WjTSt4lEU7Jo8/QCklxvEDnB0I5w18VjnXpa9RIPxJ370cmGCBaYDaFhw+vY
Qs0u4bvprTO+g/roD+4RhUjdY69qUqdR3BkpkkYX0qhXl5CgRBOjVsRYoSzBvxYYmRMTRJeOQ1GR
stYq8fIQU2uPwQ0ArlxGn5gkQGv9EG7iqiqZN72rnHzrjlNemIlm8qpt/VmWa9wY4ngJbDKe4GA+
jWSQHKDjo2CeUAvaV+DF9AfmFRpMHLqfBEI36NyRU/egp7SsEIQAoCT34RNyJ0x3/oGu3W8SFxNp
rkDsBHe0cXVw2fqAjtvxunu8baIf25IQXxgrXiyIkzek/cajPsoqpBN039G+HydlzYVtQmFj7xIJ
cbnP7Qi6GtCkgqb2xQTzUq3cI3hoFJ+V9WuJFd3K9SHXevumC3PQFK7wjF8yhnzrgDdVa48elMzS
INfgDIvOJBcg3RjrpJ6iX0gLSgHt/MRKmMExgEFUrsI358Ql65hwE0wHDHfAzV6DVueJcIck/QYh
hufm4BTevXCyFWTMheGTOIxeLYOqYBVBsQ2q+qXD0/I6edhNp1MEw11wFXnuuRB66gllXlLmUaPI
jME10Zaanw6L7DKAlxD9XMyO4ksqS8yJECcIeAmgi2YNcqVuCOo9t6lPp7apQC5WLrsPRm2GEilC
QcnehY5miAqzQj6Ljp2TlQsQEZoLUxuXU604lxrEOWQ2PgDNtWItFPNV4X1TYwEEGAD7OAwqs0EE
R3sRCb6LXavmFw3I+TQiMJQ945OsLEm0rtDKRBgtWYdO83brn1V946iMIQak/ZLryFSI/Hgwbx9O
mc8q4Cj9j+hxc1zNZ0IvopWNiSsVi8EGM+TQT6SiOCVJyAyL95L90BpfY067kqZZ1u1C8GyNzfnB
q34cYGyikGFyKp7EztYiLUG37sErtr8320VUQwGaRVClKK3cKaVA/plFxNCnKmisi2n/JR8tvQrD
rRtb+dyicCFOw0jVk/fjldgbAEkPbGQVLEdLasjA5dlFapYVEnikrZePGEJGBxDolqmV5/2KfdOj
VIGCfjErkm3NpnNqft1VtirwNO9SCsf+rzUyMFyK06IDOHSiPMtiQUD8WaHcHCA8Uo4COsxlVq+w
8aVDANNhRm7nD70Sh1dlp5zh3lpdYsDvGf0389l/jKtBb/gBabaoLFL1OvQZibRxExlnSDL+qJP/
bqQufsWK87vccqpaEStMMdFS2yHHIqN+Lt7g22p8PAgGnajMr2HINR2XPN/81MtxLSUGFqg0fu2l
/Pr4qpyciv9KKjI9JcqybkWDy5/SiYLQ8bf7xaXIvpuyymYFhaEnXmKwmWcsK9/jJAStKhzFMoAj
RXmN1Bt8pxMUQyFCBaMPoaAi0r1Tu9a6gsHcNwD854dNX0aLzgq39MU/C2kPv4rhUeYe7eOgQygv
kEUETOASPxzQn3PPO66zAMltEoLdIhIIdh4tF/GdbVShSKSX7prBPd7oIzymP7EeS6LZY1u4oWU2
OTTm5RQMFsVYPSKk8ou0R1+aUVl000tq/jP16pidamW9C3705XExq6T2ioEuC5uL/4eBUz8qgDUd
/5Ohh3N75kYW8uv5XkbYoZmcBsD+vM+YbPywCAN96lEI1UTee5QUN0jVzTmwT7DjTopS9wTj5yKe
NCQNOi8ic16gPMY0kTKFtg27UmnbzeIHDt5dwcqYXPzBrpISJqs9bhk2G99sNmHIrVgdCqW7O/Gr
Fl945Yzyflk7+esCYNuYMW0WlC0EUmMSLvb7VRCe6IE7Wm7onc0x9MpvLhk68pmTc+l5gHiP1tus
Brr4QTH2BMPpUxjerfc/+giVPcejM434BswQvPlF0DaAp/rqfCZwq8t5EqER3EgwsAxNs/V0oGck
AgYchRwO7R0e3tBW40XIN/RgjPYMXhRa9esyYheXBD72hkVvDcvzMir/SsTVYkVnUFmzOVJOvWI8
bz3k1A3HPCtJLD/NJ9AeNAEAFUpHxNGlieiFXqipY1ZSgqCJ+jyP5XUB0cDGpgrIOgMD/xUGRKNY
z5LNwLz6WrCoMIyXG1Xq6LUBnZWWnpk3JWu79feFvqCAt4c+Oz9mC+giGZJNPmbwTkE0f9ACpL2J
csSGwFGZs/QeoCh2CfhpTa6MTjKfAG2BHKRp0ea4D069eRk6gWOEZH74cE758bEPqKN5kQvUmYnL
wjev9O5tM6um/fhtHXPJaidRjZUmUmESgI6e7QYjeCCrdUfXUF7KakQb1AwaNIWaUpHWfBbQiyOc
cYHtsr+VBE5HAbBT+5ahGnfprPz5fiPTWR8bALmtEoExEdracruqwNGgh/NXTzjsApyjXqMG93v5
WJgjE5tZctRCrldyGKjjgRcDPrVgjqpXVVMNl/aEp2JOXErqaqysBm+OhuAwuY8OScz5AbxZWd3G
IqDhxme/ppBnswyzhElHzOWtl5Qs8Stja32IDMcsvkXlQndJawDbMB7+0/8sHCLWBOQouvJo8UXM
9lD9O0yvOnxt4QVrgKxCBJsuEgspPIRs7NeKJu/dwA2bm63zo9vnNdaIwWyRWv+EhxnCbYbiGFxw
NVWRTFcMYVSbfFf5rXsMYyXv34gkoBw93PSUuIdFtjEY3087NSFoWiaEY3oRrM2L+viVhi5jrc/3
80TF6Z+8nKqnA7e7L2gKaVu3KsWE5a47euv8sDgEJu7lw8yriqDv4b+uQhWIlaTYCNblX6Fvr6gr
DwDY30Oj6ZFzKreTy8RZlp7eD7PkIzxt6oBd2PsQb84B8+CmmL7XRjRCAcFFq4oq7PA776y2jBXl
75SHl2cOKSwmOoOaZMg0mM26+75D1Qrg5CEQxaIZmSdKnInb5IxIfGVvT+Y0TJKGXXbPIqAQ0RWR
UU8YFpDwelPS5rHXind3yE9Ontm77++IIp7aaK9A41LektfCOFQ+7JDCNxAHfxH/ptVPdzf70LzW
x+dj+n1LBPT3nVQVqkEnynmkPNwKjrF2nXdlKg+y+gnBibbcSlUrp3Tt+TlyKHW4EEUD5eGqQmtz
Rqoc70xjrTqL7VH06vBJRadiitBz0pY6Dub4Tr16CNtb8PafW774wgSxFSay9WaVXALpocGBmybQ
8L3EZOpXs9B8M+K/dkZGOF/dSS8lRRgr5QhM0c3CDNpGGUVcIOctEy8sOTZSJFTmS0XNa/cOx0Yv
TFuasQgAmKt6w8wyUbbMTO9qTYEMg+ccKNBFJnN7YhtbSWoROZu19qJxiVmOb4RyIVLYf9r4OKUe
BOuzMUFwudlMIUvBMTmF4KXTiMc1ECVr7dI7ISQxpihfcdIp4kN4hlbCRY1eYrO7rTtVRBQgkKDh
oRcSYtl7JhJ05IA7Yf9LNjTx82LBFtx6FBc+7P1yvrEISkrExfP/zFKy0dd0CJTybJD2GVxGhky2
KtMTDZc+XkLKuINUUYF7oUGnhM8tBgfiEMaUva+AG7V5k9Z9mrvCR52VdOQiDG6YsKqhna9kS5Za
67TrpQ/x5pNAS6gHYKj7Y+f2i6LQLY7eZX9QSJ1laVQrZaWtMdgl+KnF05ymcEFoPTqG91lmmRWk
LWDRIxfD6bPl7WhvWkai2IKWKYVn1PnZCJEz+HPgwudm6Be6chz4lC4D16sUBX/yh/C69WhLjuOv
n0Eqe5mgn7j23hQzZzQN47g8b3Phlr744Dg2wAdbGsrTrywZR5jMy/40VEDRRJVlrOajl1aF25fu
Nksywu6OoHVvhXgzmFy1/TvCP8359ltRYCH9UF14ajmWiDG9iFRDG96HkkCZBsZjajMm9L5ZhVna
xAo0kHNWDSVRA+550lgoYPdHiaX0vfrVRe4ZEF6iSrhHQ08AV636QA38T3jb0mzF+lDAfvbVLi3g
5oWxZZBG8Q1jHdTI2RnO/ePSwkiI/I67W2TCsCCNBfHJnDVUzXo1L+cIDni6rTzud8e1t9VuzISo
NqDtdabgJJTmYW8Kx1NjBRb8vdMJkZgLWpv57duceEwCALesqMAkjdhb8daj6pw+tBxczqccE2MA
iKdTWSwcfSQ22/v04XW6M43HX0NexprQ4m9Ydo4Skn/7QDXU84LDqjWYm8wwo4bvwhtPEKWluVMV
I7TbM4J1moz2Yq5a6JlbdzUfyUZQfRx6/xcofV0hMvebt/EAVvV8DUA/XCSMdiJ6NHfj3cfIIqzg
vZwScWsY0I+k5vGs5SEtd6I956RAxiYDfg3zTwdm9h6RTh/VVfoRhWvQhhis3t57GrcRZKjjdETr
4d7pLyoPtYX4v3iys/H77lrn/vK3FTYdUAhtiAf+xqq4vR7rsss4mN7SKCApemTMzWu1Fiq9WL7N
6Kh1E9xKCfkfT1addVRCwinEhRnwU97xGw9XoT2kBKpCbfDtxiavJLsaltUtqJBzmYlowFkXa5k9
qkH0L55MXNCrFy5dpd3fNl1IF+KnN9tptLo1TH+w3tnVOspvTUrblekLrUvdBTh/2h6ilNeerDSD
cvbAkX2TS8kzrtqP3vqtO4UbVuBHDMAslcEYRM75K7YTiDMjO6v8dRMI/qs/NeoR9xDP7skmkl8N
jFs5p2MSFTKf+FJObvyX+8gOt0socjRxRgV3gkG6IJvYL6kQL43cEL61PzWAycbcv8+18h7VjQD5
eVp3Z3BVzrekEx1PWjsa2YiqUxFHIXlDX2WAmzKHRFw2xPavtIzLIH6udNyK11Cl72ceRfFtCZgs
H3MKEE6mW9QX27j6QF9p9/uhMCQ0vzo/BQDQORfBLOyUcvPx5tkVnX3ehvgPopvXslRMVoXH7sfo
b7WZIiJ+Y60x9dQsigGkukbyF9o/ByuRQ4X2usBEd3t5H8flomf2voZgMg3dt5qGxa5StR1dy1jR
tu0UM0U58R/XEagt4JdM7THGgwu3odiDfXzMDwLSN3Pu+hoqnXJ/tW0/F00tG5dHzpaH7pCW1Uih
yyitBMPUDpAY9UOZoMHZgqETzkT/N/O85L8XxrtHlfLy6ccDZ8uyA8gyUDdGX6bA/oBGnJoxQ9+9
96/W2diehwUyTc3l+nYz0QEYUzd33esithol7v07xnmzeFejTBimemdJtpZ+Jz4WYu2ovjYxiSwt
DzYXLfxqPAkszavlCiesbHSw8UZIKk7cwD8ZTWSzS8J7d/XjkNbyJNLyXbweFi6WsV0yRF946kxg
4yoUl0WQgbsDA2eltZX4osNzfI1OsTu1Y+C0we87uR8y2Dm9qeCPpPGZIvxbyiVwG9nh14jdlEgR
8LigddBu+e4R7RTGibI3OkST4lERk2zoMIZkaIkDWd//knQcWRhqvjfon+13J3GFzK+dbIKXMQC8
z2fUt8X2KUIP7DVomlskrwfdGb4pHYKFRV5wCmK6d5gZ4Akua097AER6fU6oF03/2W71Ot5CPiis
wvnTLpHrT7H1PW5J/3JZyuVnudVrh4C9HQl2K/e0/V+wVhh0ATLKswEbde2pz42tKgwVJpkA/Isw
7FNVBcCLFJFTQNWjvlGgIq8fTUctF1R6pEp6KlciNPElqsLtACCdyFbxS16kIJqsP/jOgBvB5ym8
IcVtOleU+sZsyJPIUV17iUT62moOAuR6UeMWw/YjEDroBF+QUc9A2CMIoSThok9qCD09WumCNViP
drDR6vJqNhTsyGX+cB7FFv63BM9ptBzjgLyIrRgjkp1l5I7O81rXpKLGk/rI/LGd2Bew7WwEf8rV
NWrNMAoGkpZnQOlNT8qUFhOdA4jLA1gc22A/u0QoYNcJB1WRkOtt7ZjdBnzQYqHG8QmxVD06rg9s
+XineepMfzg9LiMPONQAxC42shQKkfBfwAk/2HkZXQa178uyol+PZxkXriyiwp2e//MBNvUC9BmD
nkrMk6lU+DusNN/Oxd50EcqU5eWYJCRw5+y5oskMUdiGFuqTIMYgt02dio+jwxWRkgYE5BBDmBBV
LNDX0GcshFns4BMtlVNLuq7xvByP6JHAf6+Dad4py+539yvmkPdeXDrQA0szu0ZTrkNWMkckPfTf
NEtrLgp3nejqL4JlXmcGtJ1SwsMFq3xAJ6wMjGv/gDkUB45AfqvUMunSYx/OZiOnrp+oyoNF4lmb
6NshJ/iK/IcK0PgIe8ayF5YPXLXAhhD7ecy8VpPxM/bUE0cVYIUIZ5r7oYzR87Mw/Ell6ZoBeXmR
P8jnD7Yy2p9KpTsWk7KeBTKN32NROCBVgJwElSneSmnrJ+0HZLnynSNlFr9ADOENG/qCgg+zd0Y+
jN735bxhuaCVDAADoxNh/k3td96Cq/hxZLke/lLvnlDjnqzMhbFLf1tmyDLllnmmcOWN5Xxu1kNj
4YhuhEEU66i3hFeYaptPmnQzaMZbSFU6l8T/XW7L0DD2UcnoImelUAzenxsw5DZD6hYDe3MokEpt
ER2QzK9Zwd49oZCkSe3x29CWr3R4mSbFe70TlxfuHy1lPZ4+n0cORREiHVc5aCSQ92YRkTu7HR75
55TJ7etNox8+tj5e9f9pVDwiV14adeuGrES5MsUdpNycD8jMuEGizsQNozLC06bneW9LOYidqo0N
T46PF0iO7gW3OXNLOw6l931fuA/G0S7RbCkeizG19cLEXJv1BAYu86GnVByo4V70S6CuRa5HkAbu
kySeZT6QNc5HDQfdLWaew/jTuzfIAjYrZzrLa/FPc0m5rGJZbTSuXJxoZLHiEB9vBFLeiV++hkh1
dyc0v/UR3i36HSa2bccn+T/pnuROplAomPwCuKNdx4uXLKt96kKziBBuSqh9iHOYIQOuAdDKeCLQ
3lkqUVLuRuArbHBBAgfQ4Rp5voAeedRIGPpyYo/S1KnJv04KkEPiQeYpaSP+ev3gknhK3HPCEz9r
/DbFIeQMq+fiF/ntwugMbMS/4I29SjIrnzpXd0VLsXE6LpGzghyx+3M71mtMAh/IKoV6vRN7PY0P
txkYgtCSS6oLbWmTzkzwMoPJY/TmAD7qiYnIhEARlj3HC2EnXl4jWC/mZIFfI9ma1UrdUdzC6nLP
G/AxM8Pw47qs1CkhhN2zbqc/eFaR6cyAcKHwbGEBDgJH11WpnqCxCNuxkt79dBOStKD4kBuTNllH
5Rg+7/IKxj3CS8cGys4cjLI0ao0jPTFVjA+1aulhiz3xBiABXAM8PjNhsTORUAjpRJ1+VV9RZ15Q
uczJIhP7K9nPvq5yzeW/X+zggYnoN3Ce3xkasKLkFrhNKoxZOrFU23WcmcBR9HwsoX1Jhet5kX8Q
0eL5W3PX149yvHoj3UHkmV80x/HJqL3NmtdOIPA6yJ/pdqkhGuzJj6/EAZDy/DjrSFUzS7Q/qe5v
eIb9RT6vDuXhVJbH6f15KclFvFS9U58kK4bosoa7zaPYVfMQrkJHQ/pkQ+icydIy3FfRN9lSpR1u
O17KvgE45gXn/psRxaBydDw1eedOy5VIpSscbVjFopcHRaaqh0c8r2hcyHvbQt+5XPYYuxDCFDal
z5XhUJhJXYN8HshTUMp/2En39qO+A9BHalQArn8ruDWn0eTV5pRU6LaeaFc5CzXrXqJiO2MrMVP3
/Kj1cO2zfDNUU5NTAJKxQOUvSporOEai9rC0lKuKP0S6lCpj6U7qkJ1e5lN1VnhHqzA2ab41a1u5
McCvaeZ9jh+wCrnZXKvr5saaQ2Qw3xJXC44K3nSTJxcIrpr97Bue7+qpWMMaFcPONdNnRDNvCHju
pciFB0104EePnVT5jn8U+2EUAeq5PttIpK2IrXrGlaIBu6VIih6OduSQA8oANdIFpfK7zxZZKsYu
tN2i1Znidwd432kofsEP1N6rddkP1og+ij7Oe1sA5ONqfLfTfQ9jLz/RoeA/aiUSdQp/j/lf2R4u
mLz7FPyRGlHoayDwGGuA2lmRPTbF0Bwjju0RJzC4u9UpD/FXSn/19REbcQlWhPoirc+5e9GndMva
WyS/JTd3R7E/Gfk1qxI6qQkYzSamumWaqIxGnQLkKB5TAsDppVEipTdPAZfI+/3PoVRHNs7hNgl8
ZZ1vqCZX9yihajO/loRc2r/R0D8Xij3H5yLsSU7WT7rNq4nmQiehwi2eo3EX4+WY8zOUTy+76Eo7
Q6C08NK5u6C7E/iiAaa/s4Nv/CV3QrrBrLoUOJIvC+W/P4xTDE76hdKWo1NYoDWssHVDY66y+Ctr
g6yqsnY8iRd5CR5XdnDP2PVl6Ui9L/lBinFU2U4fk88blk6c+w50PfUQPOrXugsu+gv9tA6hGz73
/+pRzHYtcMt8ODR5O7OaSo8PubGrGjlPLwQpXjyv2AaUjZl+XQbkgzN8PCz7z4Tsa4G7XyUttyQ2
nFUKnmEInWb6LCfp/ezvaeA/5T+HFG7N4Lgyjl2zcwtUD/U28Yp7ZPCtck3a3JonWsVODHgEPuqA
ZHM5hTdHUnFcJinc0K/kjk9sOTIF/I12+nmWdEpLG+JanCkAhWqQ1Z5vOkJ6iBBaMGMx+/ItuEhb
AvceWjdz8eS4lf7sN0FQNilSwqvUuN3C4H8xD4jxSJeTDx2n1hOzTDZytJMwshfzEIqWVB61n5F0
3KIt44AAEFoKko8lz3oTP3M+43mCHygzCdTYiE11HFcmC3ZVC/j8eF5Ypd8E6ZyojWvzjpNmTs/e
6MZzX6QidpnO4pzdX0PE4UKGtRE5MEkzM+1e+VY20O/HeDF2nu2xy9recQS4Pd3HQxzK3Su3vMYn
YJ0w8rAuCO2aR1IxSwnJCP/dT5ga4T5/Aoxe7Rbt8WlZELCerig9bt+vcvO0DRakdgxJxtytLJCG
hOSYbZ9HmWcMeLjdR6XlQ1ibsd4+9YxeEqr49eWvmDPoE7jyxuju1A/zJuI3hnfcsZOe3Jzn0+vy
VldN50YqfqBVszafMNJYh8HB+dK2N8QmXytFXp59fIvGufWAvefM9nj9lwoUFAvGX8GwMl421UTl
LmqBzLtEGwFfypRptqr/NPp3/9P8ZOQzXGfGoZFNJ8uPNNg16uugw4zTY2aepsbRn4wXHlnjjBmT
cTQWdp7em2Fth99eDXdOJ5EWS+NQ3bObeCxHzo6C9l+1/ivYgaAvJn4wniDnwRhJzcw4Jp7qUwQa
JpeIlbTxckH5WC0g4rMqnOos3TrnThUtW5huvL8LWeSxx5U0IxxF4vYzzDPmXjNJPldNnJ/zlUOx
WbVDMnqxjecDJ8Couh77+3+e2YL40XrfoOoIIUcLoFioxKOFw0ZRnKkpGExo/Ifrmq+THCLGaTEd
7MC6zZFiHAHl9KlUFVCzcz4hvAwVjUHcUVK6fJi+FPysDv4nh2uWed4ebUw6kgKHgbN2X9sXKDXv
tHUML/dAkD8COudrspjSEUVu3NHIPimBiwXdXMMRZw1GOAjfnLMnXncFyl9ywvwrBdNOaSBP67yw
OeZ2pueVw4aZE887D6QlE0SiDSYW29UMFbW18Yo/VBpspH8qr0nHN95B9frgQ32+SxR0T+O34Wax
67plEDU03ZGyH2wnKZ4cH2PG86sIdi7H9tnKKhegpFdfyQLhN/zG2KntPFhbfb5AhrPvvfTzueUa
k6Xil8QkDx1r1mDqUyLbd8uTHHaXd6H2ROXOK45VKm1HzXHOvBqCy42wYT4qoNIiRH/PrqVpYuGl
tK/nDLG+NEo5rohYXmIpYyzzy64xQjbnuFM2IdTTHvfeg2E718H74e6HNvD7ZHbpTNPd4kyTJmSC
LP1Nr40fj/8C5PYk/KlAI9fg9jfM07KDQZ43dv/xQ2YqxkbX6w3Z4eREdMQpBRAli/feOC2WuF+5
oxRwuxe47gqvn4oHZYpuKRx+YxS/ydYzcrvj5n62LTR0f+BBye0SvOglvyM/+u6Sb+nDg2ebPwqs
+pTh6QfHAC/yvMA8LX/H2YXf01BEn159fACQ6OUj7ss9EE3X9+IXcrGXDg9fz/VzhLHoAGCK9hh4
esO9heK7izFW08zWRm9bDtofxzNbDYpPCa03LoS6yAtkyS9ARaWBfEYxu8Z31+w7I5dthjIvShuE
wpe5VCMm07jqw57vWy+SgPIwNcMF/SSeJm23mKuPtvf9f+xFvD7dErgO8HPJWpFXAghmNapdAE7a
WnrrnLvGKIOb0mUiRPVW8wVQDgKIb8f1y+I8sczhJFTJQM39aU6Sgmfv+MsTleVrg3hCDSJRhwym
NgKEykYSqmj2pT5p6WZ3RQZb3QvYNwO/ThgxGD59Qpy8TV+9I8hQJQdYFovG5+oLw/56K4OCh3Tt
6hJLcECCmWzUrucLCE3P1Tctb0xw4l5+Jdd+LN8B2Dr3OTO4DQ2iAMhaOfL3W4vkM0Fx8wPVyyIf
MBmDSyvd4oEJMhKyXWSMvoYDRG3yKCel5jOyN3bwcEjWqzoVsvey4Rgh9EzzLu8KgoRoTTsYsK/S
KeD1lPqIgLbh47hSClfnpkZRAqrn6D7FjVXhy0OjA0hvYKgRfQVrS24KWWc8w6LTg9PKn3kTdGfe
CluiU9mrQxindaicvRKPVfx+aS8ihgzz9tdThFl7guko187DSio/1mm4k2DK45iFCdDf79mW3PHW
RUeTiLxMCf9oZY8KjxxhpEEra7552IytB4rLXiroA2g5SaZSIKdruTB331rITqMtnTFXOhcidaAE
badJghVoZnLQye+I6xQXji/ZQ5zpU+4MShErmGXXG/81O4QKNpb2ACW3BxPXNuHKcdAB5IZqwUzT
U4BPeZJK+6Tkc/mi5aYqmMyye0cKR7mLv2JDaAgUjW5LpGTm7LwMk1U4K0afe9t2mIfP75d9Rp2J
yyERKb+HVAQnZGZD66C4jWVH1vMD6hlqWrOiMkOl3cGq2fR6K5Pmt1u+KiXrikUXauxUIt/Yv5dq
w2YYuDlD0SedwWK5ruptnNhbeH2Kue2YYTSZ0by9baDBGcufJtrgVQFqtKFD/2dt8rGgAx2Zv8Ds
gSm9mpCwLq6ziPhyRmuddPcd4/gb8W5D8f0EDXDFpcz52YtHZZRmrXB/F+QVGnuv64X0T6s36tTy
c9Jz8npmA1h82XJBTafwKNXe+KMopi1z55hRW8XRdUeYqC8GBZTM6FtQOmfINU5zirOGxsdnFmoN
Gyjc7XCNRF7oIqemmkVYn54pQIBqeudYlhugOZ0wRN04R+JClUSLCVnG5vSsYY3aX5yqEFF/EtX+
6SwuqPiSCZCwivs5bnHsNXQBs9VqNLi6g6gW9e3hzuO61DH2LILJ/zqJ7kkd64kyloCi6MjxfwJe
ZXDSyEzF+jRlU8OqBrj15ozChoAldNfML2a6MpKkEHxLaPa9JO+lzSyT47/PPL1TzdiGS+qBxF+z
qnHhTsgDnpi5XcYGrQpajZY6huNZaWveU2AhTUWicRlmxhybhQnVhcGoEdUIr+/nVV74zXMLmx0G
IKgN5JBVSV/Hl3hXNtQEg0k79vk9aR0oKbY/WkgJWyTXrdfIOWfYOYo/z5EUfGQAYvwnF+xFG8LX
XgP7k7LQ7T1SO/KwY0gWwXi4N5cQeQRyYe6qAUKsfRRrgh2Z0eKtMBKZL29j1EAclvbcFfRaOiOC
f3CLY/cOmK1tyvisGPXM7KVYNlo75moLKIiqlZfuO853fKOIXKgZvkkOXY+dYHg4jCHvrtSw5PZO
6PIAYPBiyfG8hymVAfKyEjhXuzbw7u4hE0t7xj0GsEr1NwiJMF0+neGKaQoFZe9GlrD6Z2H6Wnhr
kvRsE2CjpYjFd69khvGgjNkkyG+hOAY6IfgplD99GvjsPvJ3br3GETZbQ5xnNMmkTfA3fcLWP8DI
EkU5s7QtoXpQtkBAdVz5tMpQkdEECVKFwUwrUvA9fq4CiQVuEdyx2LXrkI/8PjC9qEzsQhRc+aoj
YKh8LrwPMXhyMyUoC71bWT0OvmHL+H8Z0nkmBu2uUuOk4lgAHkf47xi+ka3inJlDcSmVxwXAlmh+
w4bUeFUNlCBFPhBII6oaJSMgAzJDoAqcKxZ2lNpm/Wn05iMdlp7SScsAkQkFkzZnHNGIN2t//htx
lwhIyTqNQ4M3dhseqHL6bptbRwgxVuQ/ZDhYioAptbcHVbnX7tfEfiPeFzWdNfTabACHr1rV7eZE
3Qw8qWrCkorGL1nSBL6W7kScha9wC76NmzyqGPSTAJmujrCuY50k/t+EqdItP1O/erErFMOLws6x
5gZMgMvrzfmnvKuXRcRqEppQR1ey8iUt2bf5oG/zztFoNLdHE/r5e6GwGVcTT9JGj1NZUiPBH321
1E7oxDXWWtH7LMIW/s1wlQlJ2oSUYvr3S/w8HrK/SY3VEc2sNjk3uu1ya1fXRf6UKSdMMl4apSZl
4EAro2eq357x4HDJP6sbzY4UVGY+1M59yR+4T24ySqq7Cs5IVNFI7cYl87F7g6pcpi5LsNfCUxv5
LZWWG9ySBjb0/6B+iG0mmMWPsq+zQZi85ImrpjYiN2EjBYbaPmEqIzw/StVGhJWsrlQX+SxwiTO3
k0XGL8RRQBHhm4++DR6caPeF+4cAB221eVDyHsgDFYtcdPZZOjd0gLFtX0kBFS5kQJeVrL0MHOmw
6Fsz7AOIcm+pp3fL/tCZw5TGLJesH3oyPoaDyYjVceiMCfphS2dUwPx6+lSfwbmNeYft0MTauGUf
9T+rEnuIyJpFOfA0DmIduxz2kT4TuusNyuMH2EUb4E2CLobGXab7q9whcLQo1zbO+ysaXIgRQrvL
K6lrcTbrRZNUSr7hJ/j2kTh4idpwSWTO/fbSVBOHD6gvEHH5I8tTtRXycrN4qJHDsBWtmchhpX6n
tlKKlEvaxi7n7YaHYvbSjCQ2yO1eZWXsgk18jRKK8TOFAflFl2Yjkm4BXlatCiozTfGfEKkhSJ0v
YLwi7uR7v5l4TFqWDbhEfo/XNKidIFq92o4TibcQm58ktx7++V7UbdRzc6KXDKBQK95fGYx4uVCv
6f+gCvam9a57Jskc0CnOnW3U+gKpotAQA9JCamIUpH0JrstL3wGbjktgCGjfN/4g9aZEog4jD9tx
dqOFFeTFmyed/yOGczxxDraTtehh6du9jt9ZwkUZ9b2CbV72b+fS/XhRAOoXPckY+wXGKY9IW8uH
BoOfCtzFw0QtkJU8XXbTtDfen12+BlpyRdfEstIy7T8wUGpuFqwiyYFMV2kCvGNiRX8xn48cPIoD
DIJCNQ9/jQ6KjLzQ55ygVWMIcbWqhBepQ+Jw32VCguE7tfu70VJ1x+xNTEarbtk7cZxx0a8Zyrar
bB8AZgNCV+Yy5k3Or7hZnPXXYXw82fWWhE44dWCmmPHO1D80WShBnBtm01gxDkC5y4jCCTDDMlMS
t+RgJ0/X7jk1w6ZW2NEuDCOPwajYTS7rQNWLhn7ydUMRDaNbUOEZ7UpyWs4RJHkpZhEDbgCtlHK9
fcaZkHI4/JWg/1LDaOMg4nq5K2gmopLqgq25TOKA/fIWAU9QQ5uv6OwNYI4gzeKlfrpIbGT5RNR3
xUr/mZZXMWtB/I90mmqPYR4IdOom/pHubOYiJmFvV+x9Lof9XkCCR5MReEO5ts1w+qmf+YaCOqRf
ItlYVnzwgCLvckXTFWKIOYOjxH5FQoYt2wY5B58MIccT3jzYZIUeBn5zCPNfEfmLj2WbWpDbCgDv
oxX6a5sEnUA/GpMJcjO4Tz/1s/wG4cHCgBUVC8w8bAV8+61NABb8Q+ACHJ5an+h8yixAYbIuCAkQ
0q9bPXqsPy9yr2zMy+u4jCnGcAbtPJa/056Uxsi0SGhJ+ydIDgLvXW2CdUPpTdsunokCsA1r4gsi
OunyxP0NOwgQtfTy6FPW1V3OYHv7OSG7zk3e9px2m3gKdJPzJf70SHjXkcGifCN4wdbjfZgaiZj3
+Y6AcVFil2B/Vbb21oRwXkRnHsbfHq/HG/9Ny/S6lZhZ1izOqhcrMNeoXm10ESLTN++T9cyvqhbK
MJSHTo/8A/sya85A8Q+unowAac+qpoKZcxy8wQL/b8hcfJCbXsYQQyfCXKQUxwJ9ufkd6RZsahIr
AvEyD7TQzgTWLytBs0snFdSE31E2o/VFjHXtgsWi/pDOiTg4KIp7E21eRe6JybL9PhCHaveMRYAY
e5f8YdkzRsahRYzicfO5S9hVsMPi0+53WgZH22joMtYalr2p+Ix19w/LZq9cg/ft51xE+lxc97Jv
yJrbLCpG7F+t4PqN+/aGqP1Beay3hXLlk1BSqKulIfS6svuzVo3fvVvDoViOwMhzAF89sn1Fgw8I
I+6teDHIfWdd2PXIPXasbFIRultNKxlBOqXGiSSQjbuRzd7tAm2f/iUxc/HybAhZyY8bZGAZHOry
gAATJsuxcaDgKcNP6nb2xOOft+trSPrZXHGQnqhpPk5GLW+qPwtTvgDjSMJuVghDwGJZXnMY0uP/
/BF1L9ts9Mw1jSQ4GHsPKhdQevdPpn93Y42OMpDywGcXuB9jpcYNfDssXumVkzRRC+YzbHSzAzbV
PJrUkwxa4PbTWFFr0Br9UXbtzkyIf/mohfgJUM87dbbPwv7+aLdwKiaZpGe+U/uyI0accTNTTOj3
EsAgT4kHyq45DpJeMdD4k3L8QNNzsdyE15DiGewDEb/xXJMw05CaMErUyraSH/O+lg9sMQ9Wq02r
dKruwHyBLZz/9+w66E6mnhyd8e1yvt4s0sNcQ2xkndOMX8uaAPnnv5A9PbH6CTwEv9q6fUFAo7vp
1S646+5+6OhpGR2dqeYykcX+4hhwJ7FjbUqFtN/LU5VlYj5dnrqXSKkxmNMRX7uTFnUSXru66Mtg
6dkV2Tmm41b7u/FlgT6Ob3mpwhTKlo3kN78LS5GMxU8ukr40Elna5/V1nB+1gIBczHES68qP3yta
RBQePCo1FYNzlYcr+EOSo9n0E0wJtPn2+pW3ARdLbyBLgy4x27Kc764TQwhYQcRCfpm/XIauaOHo
JPB88WaoY/A1+x/UZpKT3mbOJNrLAhzUnU86DX8lzdssW5npA5ZV66MDR37Kb99mYUizsvd/yACL
I9bPmgYNpB2ZI8COMgV5IBlOqig7H53WC6rH947NKCHQlRb96wF2kZSCiy2bVpTov0cAqgxHcets
ZFAXPD6LM/4hCAIyyF6JvkKgMXwIXYekUFmgWH3fGeVD72xSsXYLaHripsIJVj3Ykmt0fzENGaLS
FR5BDpCXSASg8XKaN+6ytoIegc/VaMG4Wsp0Z8nRz/gvM6MSBdtZh8UthKtZqRiEVeLMz1TiLBpF
qu3hRboJRjH8ZnM33Yepr+S+8GLN+wPWlSeYRhhH5C+gYtdvSXFdB7EiJVo5yvb2zHd192eHHPQI
UU/ThQ4yf88DauoxIFh7nVy/j1EG622V3+fbCXeRDxoqS5x+WzdX2tCY7+H3HDbMW5SwoVHaowxP
eH8VmwspFCdqVryAQNLpidvrxRzEhV5sQlBoxkMN9DMu8ipMAmiKSPQw1T9O4Ptg6vmUQOiTIHTO
pETD8VIJYpPvMq56sHlsMmDkoAK1XoQiCUo09qIQ3PBeJryzEIWv+by98RD00zZh94sg/cDUW/J7
QBp/bjOTXz9Ky3f9TdFGqyYjl0xAdPcu5YHspz9XAytXflzqdy845aAMMhLC8bRXUahs+9+KmtpC
tk640mShSXiPp3wWqzUa0xz4vd64VCzuPKrarxkNd8hWWAMMNzsj9/rzhvjSIbMYnpKGAvnFsJw1
uGihVzf17dRshU3eU1woQVIi0UTxrNzVnrMGix1MbrZJaBP9wkIfzA3SjFyOK0hmsBnOJ5lhIMg1
EZLUxwa4EuCzKcFh/f7YHFNuOh13pGl3LxahwD5pVfYi9ZBhnPV9DQDC6Bf/EifYAF+WY8AGV98i
CogtbF863ZgJ0O52pJkuG7TjxnR23MoKp/N35FxwUL5DNTS0LMM106XbZVN3QYr+UCNw72IYVEBV
TXroZsuYplSPIzSVYFZh/M/rvmXllJUXluTilNkaejuuOFNVbIXX7THt4SYgzYgOOX6Rsrm5cuQA
UUisJkUlPg3SiK95Z0Q4HczVuI3puICjM7JSLPuZUxeSvzK0lAwTFIGXJ9I8B8LMkDmqFAmPaVNr
odBKJSXVGY9bENq9d0U+smqwKJnrGfd1lYSXCNzHqYgaHk+PRTaM6IFk/AyJWsMuqGeQeB/zjzls
YBkPMNxJULTV7SFlc6a6fQqbVvLGRNxu2mQ9N5aDOywedukcrtUXKUrg6FaM3Ld1DASW774ejiRO
SbWu3853Q7NPML8lr9slzhR8Qnn4fw6DcT8sAdM4aEKGGwTxPOE+j5wnfZolhIXan+NqUBGxB0uy
nxll1tHor+RZ4iOO9+KjNS3Vq4eifrRPCxnaa0mVbJwc9J4e97+eEa38BBZEDX/+RiiDmjORICsh
hg5dQNtGr4HgBhXaJ/rQhMZsyJuiTugJuYsC45LjE+M7+QPW0BPcfHKasmha+nscpBDddl0+L5E3
Jcos4WRQU9D0tCPHEkhabJzttwPVveN/nyOKFNfGl5LqHQI0oO/LLmTp6ZLZtY7ErRACjNEnxSjZ
zWNbJw1MHWod5yi5cZiV1ESxBeMw4lAEuwTPfwUM2D0g4uQKmGzeLdCBiyouQHiD7RK0PKubwogW
WYhUL1kg/Zh8U/Aeaqmg0DNOGqiG57NDP4kaHusuBUmIieejJPcE8hQwPLO6/nXpX38+KYo+GVAE
IBxFaWo0c3/Iut4x9E1dmAXOswDLD1G5obn/hjIaxz2Ue7z8sq83lWZ0zPLjJ9ImWI9SYG4egiGI
Ul8s4GIxMR4R6QBX/r82ERzI121LwkacarHEQdnbfasD6Wv8EOa967Wh7YjeYE445GN7n66f/hOB
2CyvPD/MhmKy4wASoywO7yBh2qMl2p6gpYLPPuZ8R4uyYB2q0bMrJRgZhR7KMHlCAarGgbwyt1ol
p9/vIx8Nf/xpMYjPJFl/t3fyronK3N6SeztAOZtykrmrnz4vm6UWCqQL/VR8f2Au/oi9F4cFczLT
hQw+r16NLp/LRMprFjeLAgSngr7XtoNQzlJZdF6YZcsDhQmaV8pJdz9vE0cXSwFM7SwZJuwc1gTI
L8c6FR786v06Enh9ytcN8ckYCQ5v43QvxBKN8X5WS2lIqC2rsbNlJQW3eLfxy6uJ1uPQryLtvHRY
H230dcmxAh/+wnXH0ZhTMfNttaqj67Uo+JGkRRxRA2MIvfyyAtzfhvHczGqgNUYvHy32SVorekiq
aeTogRbkwTpuMEH8stzUqq1CSlkGf4MK2ByViBUdPQvDGO8gwiEW1W8x6HOdY3VRzXnmxGT9wErL
1TfRe+Mj1X8WCzDGcbVuv7LZEpXLajXdfdIdbbnytErgvZ7M+Xl4nsEUV4KXY7bSfsV9/wVQe/hH
KKXywaX3l7dGiAuJ1Z4QOkQNNg4qB02OJeQEqeqrc5poyakALbA/8Gtq4JFX1nYCFlRVVS6fwPgM
8Mxj6988tVVLAvscPKpD5IZ2Px47//YacE4D3H1wsjEAFw0OMtM3ixkIo+21UfUi76my9s8IkbZa
Bd4HWQbmTpaSVJO0FH9/fCpdRGcXdGnOXJbGWDIcxio31/m9PEOqFRJsBRPOvolql8ihWl35qxqo
0wDZnhVuOR/IlGFahXPhgKBHyIU8mPVuWbMQj7W/c5kHqmmi/TTY9O3p1ROCk5+V/n4bqJx/faFa
YkKlrNwYJiu/gpQzp490eYxa/44Ui3jmRceMn6TkKxRCJnyDMlQLel8hfgeM0nKsGqcLOdKdkm8b
ghDJsEytsh81f43ggvS+QueBnA+TUR5lLYBLfsWf2AlIBCxUSOg01KpUX+D0eX3Pqx0XFcqqrwEn
8l4O7Ci2tcXAWvI2S3jVgLI474HQZcruIjRR6MdgpeG+j0qxO9hYTiMSXnWZwDKfrSalsmukYLd5
K8BJ5IxH4WWH0OV4UIyC57Zwp+3X2C//8usPG8UJDhDUrYJ6VZu1mx5rraw3wYscQbTFz+aaHwz7
TluFHFReRVdo+5+791EbIiRL6M/XC0TTSOsnyPZOgcuT3elJ8fXt8ay+GDZWLOzpaXpGp+X5S/NC
OdMCqrQa2Lx6oYw83mEGqneLjCbkaIMyQiiUaRehGmfYI/qNevPIwXDhuCZ8LnGnOyWt4fXtOumq
XgAJ0ZgV/fm8m9G2HFZaCsQU7xox9yzn1z0A4iDT2uxat6bnkWEOUkVMLdrFCpQwBhk6fFqZuOVo
ReBx/CCzwLOPbnC4QuJ0l8FvUEhlaxGam8XGo7Uvyc39ZI7Egp2bcEqwQqIQAs1EX30XdesheT+J
BHw1kw1i160dJ6th7Wwqpo6cvDcgXhwQ/SRzUG5/H5KUaiUSmLp9rJWlw3EuyH8pOyyIyyvAIiB1
RdqLfkf4uIuCUbp43rOrpBTpojpPoshNwo4L1wHuq7KWPyKMYFyC+kr1DhYwY0ay7Ym0zoJ9QBSW
OFVzasCgMGJcwA2bqRuEuzBSjVE4su1JUocXhQiFQtS6env0LWg81f3Bg6wY9px1Tnrw/cApG9rs
4U13MLi0ZaWavE4lqiaB4rpjzoshujwI3Ui2FuURfRW652mI8j4fqIX4kmPoVT3BLfNPsoWtiAtV
Z1vEnuj+qanm8DDe7V9lgTzXfa5oi55zMUMILvf2qjHmpcbFvXyFKS7LOBpUH1KQuUgM0qWNRVm3
mgp+7MGzweLyJs8mz3SOrkox0qZysAI2Vh4htwSZeGafPLeq/426GpwHTtF2QqB5kd6IHJw80Puo
iJMyJ/7cpigZ5V6YI3ZwItkn9STYVCKO2qSrQPFPSfRbgKX9ryvtucj6V4MTn1csfTenvwc1atOO
rRwWJWtg+5bQQOsvH2dGHN3L32yXUeL9Ua/UE5Ok1ZdXFn8EspAueot2lqo5a3jTFuEQYEGezk5Q
tINz0OKAojBCHXW+bVgEEWvkjOWIAvdqrTvLXq7EcuFfFQ01eBxOMl3LyMgnjtSBPDU3X/JkSHaQ
+C1053D0+eiZD/jUkWPTW62LxlGmt60aYE73RGVZvyWuFVJF2pnVxcB7+ouMlPL6uJkPJhh16Z+g
6moroaFYNv+4bh/AUi4eDQbJDAWRJ3lGzatzEoirpqx26ic3lH/MRLF4I4lrGnAQtk2l7dlavgwt
0RsR0GB2nc27gcK1gROOA//j3aoFJ3ehwF9G0BuPaym1yAKu6rlkYej/Wm2SbazSVl3zpG8BQeBa
IICNjpR1wTytiHCL/6Pjdk6LIWl05m3IT1jHxe8oCc7vhIXfOyKlhOsIzLGD6Ki9ayT8kDm6IxZJ
162XN6V+JHEFihXe2TNRs3kEsUqqQJIp2JqQwpWUcXx8MXqh2mEWZVVdaqxpfEcLoJz6xr5+ESfT
mRg6y7n/HSlrhHaWlPf9MblVig+GRVsbKNhcLRVdAMvB1NChF0QFQvdN+TVyQnYPz3AAo7W6NcTw
pawoj2R2EgdLEqqr+BtaTxYpqVl8pFw9m0fxitcsu+OmdAdluuSxJGW5Iolw6+/BdIw4TC8KDmwO
aSXwNOt+TCsZtyLim0+OjNhMfp+4JLYmW1Rxo4HHaJBNynZEd3gVNxaDi55sJUjziZPeKWBXdWpR
ja/YY7DSg/kCKntHPQkKjfSHPtFe5lKXrGs5tir0+3OyiYlVfShZtKn4yK8z9vESbxlmhj336R3C
AZx2Ao/vdOHEg2PnCYrG5Zn8Bl8gpX98cdnk3RqXi6JIxuI8SWe172unJObcIwY0Qo4OYqrr2e9S
nVRyGfKosTAXe3eHOtg/jLKd0tLF3iZz8GU2xU8WxxsWCzUJTIAaOfed1YgC5nkniMn0GSwOM8Lc
0W6GNl69zE1Ho5aTKqGawLqhgFo4ODWd4BLf1rC4ETrVeSCKn1L6OEr2THIIDj/uPjPLM11NpokM
fZcqjRJjWFPaBJImXGiDVTVDyKJaVKHuOwKs0PKvSDapZRwP55LpfbuZX9TSa5B6ODno6gDjZB2s
+3s2z7vKhcOdoCu9sk1G9sap5+lAQcblGFEDB+FSqluQC7RBG6FUw1H+KFpsXLm9ddoIfdSpA6EP
kRHu0jdpmuuhni62qQGp0XaDpZOXEEXRQSmZzmoe4Z22cBRKLZZwnl48m8Q8+N/8/gPin7l77FcD
G44bYs/XahqJOMg1qs6peADz4lXwp4DnTd6d7ZmpxHmiTQ5dU992HJOVnA5BIiAYF+/NA+v7qtwp
PN/s56KRKAlqOguh1pNZB5KJOuaLMC54N/nPFvUjpC+rM9cn+voXQ8vE/BRissbjAlIUKqUchv2x
mdfn/POBPrJ6t36WeIo/06vdGUDIjXbo9zawP9XZaO6dLC2T0q539f5GNEZ9wmqPn/7/XcD1sYOG
0udtYuq4ZJZJ5wTlaD1RJq7IWGClX/tBRrf3pHDonvX0+mlOR1SuxeGrttgrKAcfLzYXCsLVQ108
qtpLinYBXDhc6pT+fWmoBt0lrcfGOap5/N1kWXC1hVPROUjdGCG5cD0kP89GiK/EdMqhjaMpdE4p
UWRxXxfYnzuAJcm3WddaGfBaHmW5LDrCTsEBRllGKLbvpgKbdBCs8QbDsRSu8UoZaHrzxpFEynY8
cWKoriObT7moQPQ1hJhSX7fjIH6M2uwm3MtCCTeM3MwdL+QODpo7yXZiAuGnLmw6vgCKkGUuQUKd
LwjvgzmNgTccZTuJDXEp1tCq57quNEdUoVVlk8UkcdTrKZ68Ve+WjQgA5g1pF4miG3V3796Qvolm
Suruhb93QfDaAP2UR9kqNWaWP8+XaizFPk3s5pmylPKm8sgFIgCBgsmIPGZyoHrPtdA9z3M+A4qQ
d7EK+s9Ee7PZbxEXQ/7O6MWMopbUMEGh0q3ldQPtc6LTjFzjE6UqoT5VAQZvPU/j557nlMi4+sdM
CfAlVym3JDx7eBySNriqVCBIXXthMCFOnyiiPAmo34oFF7xOmWhmf37J3nbIVIShUOrss+d9Ueb7
c+ZDTrHeBmnp9cH9vHZUfG1HYSqr27Y6Vh4jH1uGw6g/ElleZXB86IBFYxmUExeR/U2RtWh8e1r6
n/wht0NtoX3R+KQiP139g8reyJZUHrrd8nMglClIDlDGQtq+2mn1Ht5fRYP8oWgrf/x+4LyeY71i
yr3Oyzk5nE9SstNjjU4jIhgbR+YM9J6BYbTinZrBf8Jn5rsCANJqLK1Ib+zw3eA8RfbU/wT+TO9v
4QmHkFKFJ69ZP4ajH0ox0KIxdgaUwQawN9DvJ08/8LRb9xH/kAO9uydetrMBO5MrcMO9HXjllHam
Z0tZxcBTy7ZTGsEXurFNYjuOAKi+DAhHNX9amhG3r0P8WmcQbDGWayeADMuiCfrBFppr0/C6DBrl
iiPRySruwgCWHb/BETxNyko+CXYrZZv5ehmKxMmX4KuZ/g1bo/vPsXfv+zoa53TIfxEzMIoiGMD2
zbTA66bTdjGmT8I6IgSCEGoXui7oXIERAMdD2yhUvG8qM92JEM6Ysmx16OGwa/1lGefXodd3192p
lKQWkvHf3XxiVw2H8x16iuIDlt77fuu+8qHuV25Pe687iuAIyt0KKtcAIjetFjA87PTBS5H1AdLe
AUtEsqKFLjQBcdDeLvMMLaZgqgXy0vH07etjPidKs6w89w15xhN2rSe0jI/yCd/qBW3aDTvlAIEj
+0FsFq931yyko4fUdsi/IWYEWFneuBDoccBZJtEBXFmjqCkXmh4KaYFZXSE4Dm04Hm3efEiozEFW
QdHLGsxrbsm77BmQShHQnifs3w/oTyCcd4NVxc7dA8oUKmGL+muUeYWUwiSBNLPu6xFyr9vK0wDX
iY6YZMGwoa8eqjION1J9zuPQTZKwXEUlhTEsweUsLStU6HJrrBWrsGBv3CY1lDD11x14FSQTNzC0
i8tWtAiBq1/UwDAUa8OqDb8Kq706jJXAjkL+ohBGV3tjssKoXG40MOP9WtImlaboRNTyold+bvaY
iRgx2t/8JyDY4QJSkP1M1zYfEcudl/Jevltp5xamguCPZI94pK44LVAlBYSmLa1ELeMNJP+ggM3n
7QEi5f3vlSXE2ZJ+PBkUK91sDEfHnRCYmJfje3CmgxVu0mneiryi5kfLsX9BWfa6mJk82z0I5ccb
veYcfccSPKBGxwxZyq8pi9/Rn1nHZ0tvytn80wXE2tQJn/dQYZccXZKeScNDat2Ho9JXyus/VNOt
h3xBy3IJxKn79woQ+S0T99XZmhihIEXW5D3kq87w2VGULAmbN3+73ijziR/oFLN0SkMabnUK84gC
U2EqyUW/tyb1UlChFqhblCY/lSNSOpvaGVRfl9cLHiWNY5Ji1eBGoEfkXOp/SQaucF/m6Eow3PHv
O/Mt0X/4s6KkpiPZ4h/Ok0SLizBkO1ZDcPrzfUEUHlwrBCH0m0Vs+OXx3d+y0oyPFFFALVxW2jlt
Mo9F/YzmRerSW9LnKs9p5GdQeLMh3453Vfhom+aLJJdeilm59ES/HmOgsN1D26AAO6T64MXyRbrg
xHqBpTucGiNmsuWK2Wg7867fWcUMA7yDvbzB1PFsflQRXbGEX5MO21zVuJGjwJ6T3NCJQejcbtyA
bjEo+sOt0LmQbTpYQXyK9c/UEqWftEra4ND/UiUpnhwZP76Zgam0yTDCFyp+Zxw2D0sR2UnoLC5Z
UIyUxuSP+kkbRxA9IW4acbqwVpMprHt81hOVnOcMQbwZ06hzNiSlW7pTGT5a5bUNmBH3aIiRo3z6
3DoSkoS9166HzH6FFN1RLcgqKV25Xdgu6a2z9bf6YHsS2xsyfTWRk2BZuZBpOFENIyZtAucDhmBQ
7btIUdZ0rRcoNVcwDRdOTwBZBVewK5gRCu6K9ElPpRvQ5KOSbQA9gMzeDuyMuZ42g5Y55lOk74EN
nHm5Df5ImWKUoiXVQkrbeboZmFKtlNV/ESlk1kZAp97j1TTNXU532/acJ4Xfw2erYAv0W5/5JGym
B46z2LsQRe4ND8PtIa0XrDZOW2Yr0oEXpssfa60rpvlczj2mvvWkgC1BznzNXH4mUhQFF2HHePaI
YvB38cu9yghy3lalinaotDZ5FT3U7VFEZhE7AmlOh/E0zLTpTaMRRRa5cQpDpyZPzHebwQriFdf6
y8n0zt+ElEII19+c1nAEtHu3BWSelBi01l+oyYGUrm9oIN1fZogcereKMbiaacQyA8zM/JqFIgJQ
+O2XgNr/RUIODALhkLc8d6i75jXkQUlHunKkZFwkn1cFFyOMZx2zvrBGYmeRiYyaUz819T0ORfoq
E//SeMpLyDn/KdDYfuMDQKhhNG+ZVjYoM1bQW+KSxkuUy/5rm4ZzmE76WX//S4XHwCuHAIaOsR7r
JblyAGhG4uSrboudN/clAJaKZCJ9DUSSIjz8BukBnQYyZn4GihNbkpDKXVMVInNURrujqTjeWZ0g
aKvuav8WllDQA6xOMaw8a6093cTwcbAJVj/WSZROVDf/2sdsd20ai7emdW6XY49QJFtN90gOFoqy
HDgTVAn6+mnLi3ti25MXqMd0wrHRiM7gnwbA4tr2cosGdta+qA5XBarxabS1SxtD7R/BaLRytiW8
r/+5GSZ0DVY8mpe01WTxKoNc1hPsMp0Fh1eT/xV7+Rt/sxsKEKSA0m5egRn06L2+J8PHvoziCYcn
urSA80bJiEfRpH7HuC6s6dgEe4aXzoI9E9rrykFSUg5caKqd07BjcKsvPAwHb5uXNT5GHghFwSAg
RIH6dlkxoQrq+2j+nlDLixv4staGUx6u7wQpy1LlgI9kwy4w8vRd5hSw/wInVPuTh2E0UH4efSLs
n0W2fmXxR4uAeJX3/PVqirZmyAAujENNwn0d/4K8w8j/vwxswsZ6m5tlq0mntYChzlam096pNdsh
riddubDq9mUo67/8PI9cOO6P8c+PNhqwpLv4esJ/PW5+KS43m0m+wwYC/DJml9PMA4GrNAclVpJ+
1HtbSjfx/bTaWBxkrwzSkm2abzS+nojF/0upcxsWzaQJl7inuOcYitqP96bP3zx2LEAwdq/KHzsN
lrsNy/oPjLmGoDwIIln+hIjiHpN4zAkPhjxJX0e0hZQc4lXIVNL5I1Hzw4DNG//hu6LqSKOJK7An
7KjARAVpiyYj9vfh76f+DALaS+9DPoBIbO3p+noiv8x+fqjcbLg9Rhs9y2vKm3w55OQny7Y1rEdO
H+JBnd/rfoQdKLYMRJJpDfDGzFcdbKGcqop053xS+/hhSXdKxPo7JhP2/B9iHzV0ZJKiUcyxAeoO
oR5PVYchizwDtHW0SXS4bz3DZ8ui85vT72Wcckq9Xb4jE2zqpTKwocOSzzCuQ6p1FE8wq8f5DOAy
E9VGqGWsqmhxou4xt8A8i+4AWwX3qGqGOnNHi/g2JN85ESdk7rZqgyciVzB+eOqefXF/EsMvJwO1
lnyGyub/jpUruuLW0+b67a6lq16PWVNLrciO1SBcxz/HzxUPzgpzbrpefFnKK/DrThMO2BtEC1XH
zNWhRd9fvf2egbWAyTacsLq9V+FHn8T2QFRBOxCGuCSJ01SrnMYReFWE18D3RRCftT6hdjdf5s82
51VPRwrHXMa8KzTYXpiiUYr7j5QQbLW37Fh4mg62JUrK3pdFKKXvLtwqDBeXGS3gMfOqaHGF6WQM
+cXLHuMqLQ3XfrUWlM32EH6No6LJ0TpqS5DDuZgvsGN15+OMTj68JBwQI/81X7SHj4L0k0MUoyUh
nBhZ/K7MB3qFsoKbeZTILw+QWHxcAPUtXOMk9eIFHw9dp4GXfc7TrPCTJfe4twCTb1gaba4Xj21M
8sz8UdqjBpRZwAM2eDgz2Cdm8g6HZc/fWFgbM9yElJUiu4eQWWu/PTOyYstcRUxBKnRpZAYv2/Zi
N0AzJp/yIblELjMoMk/6Zl0oD6s4xPKlNUYFEOtYgNnaBy2PoCQFj2Y2iClnIdXedaT9N71FCXKE
Wug7mXgAnK8qbUAmnL7xqHNxJvQWcTNY4Y/fnBXPSenj/JKiJTSx9b3CUoJC4gz3cukrkELMTsVU
18cBgNXCgB3yjhQ7E/whPSdfzXXm18B3weDy73D4GOsaMMEU8dYNlnUhKq0kuTlrsI8V1H20hXb0
kSf/QAhoWrf7Bbj6p//FIxWfsqZz7+/1TFPZL8Te7agV1xMvmltG7CiN5eIwF04DcD1eFM8zUBU2
f5t8P3IrBudB8c9NtikUrMb1rOmGVOXb9kl3CcEctkv7lzGE0/NiJg3hlDa7aKyVTazuMht4vwHr
T8cULBWT+3T6IsSsPJA61GtGLRUFoNnbOkpDLwZ/9qzt1rOH2LatzI+GGMlZ+cX9g2KFXrwuTIgC
k4W6zobx7nmCXwXiPtMpmkdR4rL+cVcrBUQCAWoConex9JdB1CSp4gdqOA9aD3x6ctTC6X6EQwq7
UkZ6BRl9zuQM0vCV/0ubAIsOjPXa0oY7FfI+4pp3tTtu70Kxl4u1FBKP6U3caJcIBsZjtmqVrYWE
YuTqee1tDHGMR7GatQL+lT1fm6ynhkq8FRjU6TJThI+SItSeEcLowgfLwRlNX8tzkKYmEoX/yg20
cMtSD/D6rYds7F3YN9nTaQ2JsX147nRIWYlCtTMS/r3v8Rf/0nHQoxLFoIrhACyCRWdurL3qJ/mb
d2mQBTb6QTllwq3O/RP/t8LLcrinhKEEQQbuNJy/GuwXBsR+T5ygQTbMtYNJarzMZS2ilghpVYbD
GUU1jcSzen/O841qxEqL3uUWIgo/jHtySa4oWECjiYOu3JaNGL+fMr78k5o2Ve/HnMEDZZzsiC80
Jg4Jt6VZtn6r1b2COt2OlGYyYwJL4ELJhMiFfxiHJBTDmqkFzTicXZcfk/YkBpSakw2uNb24/9+a
9trefxKYicXyc8GWNB4OX4X3snavLhku5X2QdsH7WeVWpH3yriaPmVwOYODrV7MKgZXOVw77uOpW
69FeJ1+UxjXGe79C25Pafvnm9NzUlv5tiA+1k7ODg67E9nCCjNs7agdIxTKB4qr58YERG8FrK5H1
17/RpTxYTB42NhEpvnKBIe54d+En4sX8q+uVJvTyhzGOEDYFMynhbfhDpwVvnOWZwab/XQkbs0aY
+hZf2PBAP0c8WBMnwYdssgGqzRpDSsqEISdCLFpB2Vc06xz73rgVvlBsmmSvUv9zaYeSJREgJoAz
J4iZgiQmvNBgTXHOnjmc6YpbV7TBdPEN5Z9YX6yi5S/sjfR/OKl35uB70PxQKHqNngnQvWqq/cId
9PW4h2/1PUQDcAb5PQ4fjskgRBuROs+7sZ1kMMMGA/8mnnCR5M/KKTbPRDjPMchn7tnYvs3cqtOp
1YPOty/RkBdzHsjIhj6BXgWXIDeNu6pqMzWwjcEdiCDy7DmU2ATXcTFSw3H7kyTzoKYfGwqES+63
19OZC6mBTDzRVK5klfL6OUXmGekNhJ9NvpWvggAfnbLulVP6fBbnS/imIA9wD79LsKciJ6QMBf91
wVISKgUaANRvFXO1TiaBLSSkYfcnbOr3U/0ruWpxHmUeSSzXa5yA4+jaPnMkdD9Jsf5Feen1LHAD
6hxQccAbdoTf8gnIZb4s//q8tW75UqbZZqgDhQdXE/zLXPW+Ib9yTHW3NPklcju1JazDxsmy1DWw
aWyFDQaC8dAJiIc4YKXYekZ1P4g+kQ34xysN7gKiwhh4JsFhd1Azmbjwz141VZTIZXtT7JU8ItPC
igjdx8oBIRU46oPWd91Fhb0zWXHKSCQSejjJAB+iprT9cebECgt5cW9QSPP1OKhcpBVMMCvqJ/UQ
lL9MB9zbX5w0a0o5czJiARr4qSiIrSaHrp2qhNDZnpJPAgYRJVnu4mX728WUWvN4aQ5KwqGoIYgD
L95AgfypTbPAvPL/G8zfeCdsOG4wwWWAsJPFEvBQ/B9AcFF/cqtgUehuy88/pBMWX29JdUPfXzR5
Z0jGBMPRYYMX9nG0n/J4rleJj6MR6o+quXTX8BggHaZQJgbWU6LDQn63ACCY8p2rp4NCd82W2N0T
N3ZWHNR0PXGTF6y87+/P2dntbxzjamzNC5EXYJLdP46GLP/nAUv8gRA0cQlRBq28QlSDFKJncM5W
BSwSJSGecmZ65Wy18xWFOUTWRTAKWmObFyiUNHsZAeNB/vB5PkBUBrQ9HrP6JqpJiTM3/ik4/+iG
eNbj43MqER4YhicbQEjUkDf0Jbeu0SpgNsWtlD8/ULQJuC2Fgbc8H/HYmwjmT+rFkrj9u4HITBSO
yYF80LfbZgUMegvXJtfuGwfjEvfCh3i5wjXxJrA0HsAJAd7/QClAOQ/ZMBycMBHI7P3ipJYWhbFJ
h2LAQlbPTJc7UQF7FTYEcsgfWH8eAP1WcitcwnBRpRRvt66qcXYyNi86Mbh9vndYf7EOITUaz+28
7zaemJPtmz/1SUH7SUa+1fEzsbnpF7jYQikkrWUa8pqnhZq3JX9A4946O4eb7J9kjmEezzybJ/Ca
tHdNpYunF81DkoIvVnGU8b8WCCue0GWp15C/7ZoqbJiPI6N17iZADmdaz5ajhJJhntWFtdzXi7y6
7Mi0xRERgVlxwsG2gJSnhQwQyg/oI6gLAXa/ij86NNOY7b12EFva5CqAsi1mY5ubQ+xsnKDDEy06
p4o0zfQJpNjaOImxK0OPOZPL6r8A+Ty9Z0uqrwiNHXlnxWVjKBAc+tIa8UKwHNXkQtARRC1+RW/A
SyJ0jQa9PUGTrKjbMbVqsSJFERpwnVzZ9N0YnKikTCxZ62EBYRxRlmwF1a2zPaKJeqftTDaW/6/4
FXOdlazv5lpmRFXP3fO+AhJMlrHagAY4RbuP1ZNsKaU40MRR9LbovYaH816oDZO+ks14cdDQDklf
KT+8bib+dg3bRMbCnD0b/KjE8tkOrPxv+YiIZa7/D4+aDcZK5SQW5bxDg3AzZSzFVRCGJNiFuUrR
Hl0SiONJxrGBo3ngo1GBLBDUWUhCotqlE/0zRxFqOajkLITYjZHMVTJsnr0Xnp0asveeGuEzrUV2
5WcNjK4Lo4FgaeCwLt3ODeqAIZ6TLnoQ8O1+cq9JHsp/LBOi9IDWIkcRu9glpqGlA/0cQXXJ4IOe
wWqqhv8YCwL5yB2wYnY1/QQnCm+UXdKR50LUf52SZoS/cf+mI/xRLNllKW0hELwvY57q+7ZZPDds
AqN4iZfxAhybn9hyga4kLJuWyCH5Fm5+ny+U4nvqjKdEXmk76q9f6e4HFJwYsZMGFZGS/LGmqbCP
8BJZdVHcMT2OSUP0JCsgQaBFlpDYTEBqVi/6WnUzWKKNkHWWNPlPdDrmqje4Yanl+EnA4u5H/bFn
PLbsglK5ajvMKOil0pLTzWZk4azGf92i4o52N39y/Wo3dCNY+0bB8X7Rs5JuJ1pgZjUFLuU/lR4H
1ZlRJffcECGdBsKWGFryhhRfmpRuOCR3WO+Tua2iKQC140QchADBqoKcAJD4MJqZ4iDDB50tOIRH
P/xcSuL/Cps5XnZECe0W9oUSzzbKgDPWpm0/VlAmOO9ah7k38r1ntVm66yfCFhT9Y/m21/92kLxG
NZG7I+AA7dKt+0wTfo/mu2J+4MhWQURF1gmtXoUNpObSDIXofILMfj0EJgURuXSSIydq2a+T1uC1
BJmaVnZ9nM6zQI90/ONocDGVFuegvpYvRN9BX26/35SW5SjM/Uq3ZzHU8oCFuGlkIvfa0TonC/RN
nYWCT+xNr1mhIbzMAXx8L4sBEHCkcCpC0MGSH0xctPZR0wKZWO1Y7Vunbo60pNY9Os9J2nzT5Mzp
uhIdJH+647XWMpxjl+43aXkN1hmpmvXHQngUoVCaYbeI/oAzskXgd4X4LhLSBtnDuKxRzsHYFGWg
dyyvSuexO4Vg806rgFw1ojq8x9Hrbjhfwf7eQNFeyDPzUFMwomNFmGfBHOr4Bj/NWOSd9zxKZPpL
ROansfwo1mGdnOezQDiqTLn17ylGUO4jEFT9hLNK7icUPzTqSd9tLJs+OP0tRTYuLIjKVEBZ6A8y
oBjviLRZEMtxsz2vkm73ecZtWGcTMcerQ/YlUyBJalLjQSOX4ILKCo8j3TQuG9/OOQ/r9qKeWvlA
u5V/LQXjRQTmnjCiRKY80LzPurMr5rx30ZNaOq0IAG5DtyN8Fx7MK0HwTYvc+gBjpJbLx14welRc
vONpPKms67dA3+9RTTc8sHk0xUseINBb4r5PSZQnwTxuIkuf0Evz8oZBbOx6ZBQ+mBal14anxTUU
/XPmKZ2+QZOjbqzh5s4Qas43coQnGrmo3vwUfW/2GTNkiBy/g5yf3AejUYYNXm3VseioJXc5ySQu
4hX2WHi2/0zucFg2ditK91LFhOHTwFbf1g79BB1X/mB48xw53xbzrnKRFVlRYgE83K3PyIJMsuLt
Wr8UfxYjY+dHLMkqpSduvqkw3gsYSRnuq+L25T674Z3wrQPf+Ex9BkhU4kutg5GTaM4XRJ4RXBes
QqGyNFyNCfVWFRTfmsvZKSwNG9fBe06ulBTQbVrBYkwNSejcrFOTgYP0XktZ5A7gz8miWGGBCxjY
mg+iwYkr+yux91c2KnyZMjDvaA2lMD6ZPTDgwq42tK4rLomK6dUS8bR57m0m6RoShCsSGmLhQm5e
TzlAxMDkaTUlBMZvSucjCxIChCDPPgTgqvAVxOdLtkIM1mMzQedtXT1VbBp453pC2CDSnOTFQMUi
3u+B1HbWeu18sRyOaa+40N0fa9k6yS1sFgpWneHAjK215SebXnluNNXUVqHr3ciGObwINXLYVuRS
MwcjjtsD0jKfta/sV3tqVkNZtk8N/KGTurJ6qiEESpe7uG55m07jZKBeZLs7RypaVSgsflDJ7FU1
TGw+S0fed+mgtLtPBcwmyD1f72ly84PjQBZyu8hzPm5hbQ0PUWTDpevtG01SBb1rGlmri3kpoKdN
DKJK8yzf/yMOouP4vrIAer+j0SWJfITzF5EY56ntWUPJftLr2kkksBdXUK4GaulsE9DAmxfZlZpa
WOzxkWo2AQ9YEnIRMNTybHZzc/PEStayDgKy/Kod3tAcE/WyB+yXuVNsFu4WDNZ/MLRBU0pgr8lp
4AI8XvC1FXyDa4/w7b59mpxFnK2YWCBYD1vACl2f9P1jjidJL3ZSXydq3EGyy92HYd21fx2X4aYl
PIuEszVRmBJvRhrCptcTf3tW1QGBvlTMxg9m9xWwYqQFgHCzGGnVyigiQf1S0v+8MDCuTt0Nn6ai
c7gCRLn0CJ+FaGTjsIvuLGXHT1J6PRg2exp8A0q38rbj7re6paT2Lj+08ZGdLA96wYlZt6SB/ZZM
J/stopn/3ZueYr25V4SAJYr/h4lbM6VtBHj89i8v4fD7I/lgd81Yfn7diWhdjToPhMzQEcvAHCTC
lKzg9AZzynnPdEmjGo36DauXkXtC5cc4N9yKQh0ESxWTwHq3ArEsjWtrJPrBbBk13nBvLFKiyLdE
BsVIPILcx6l0sO6DUdYIz2HvPHqPNziGJ+IKy9CszHUKpUl08Cyxas86rA5/QN3YOtT4Fb8xJvSv
Dboq6GgtLQW+mM0vLDYQJW3EmBekVhIYY7YQtTUeq7FaSkevJdxVWwVYHodHuqAbbo0473+jJf9o
p7IaEe3NTXW5UhLzMlVih/ilY38OSck+RhR4T4h+HYY/9upBT5wCj5mkKFAWpn7ipEoBJxB8y7uv
IKcKBphVPL0NTTKds5/wWuU1xKMVvHvS7VjLLb0BoisCCSFV5Rt1Lqnhxi77U0iVvQD55fOZWSFW
bh7rhknQ+yHK3vLsdRS+rtRdSGGea/rc5Z+wVcfqe2Cb4hrLiJuDl7aIUTwcTUkGiDH8cZxwrFqe
RGi7CJdm1eBhOmQ3+JxM0YWZKsx5XpevGNN/G35MK23ux5MNFoDQ9nBEoyuD+4CSnxm8QeeoXFl/
lvIqaz3C5jCVSLQ/coKv2c4IuOLTgXPXDU1wJCdeWfn1fwieBCEGrN/KTk6nMP1iAguQI911f3TB
8wIAB6S8mIAXhRm5UNFGvuQ8Ly5UNQxkPhv5Xqm2DZTiP3cmoXOjAcurxQUEqs1x2U9wa7PHtBRZ
9vq0VJ+ARmpvFI8z1XAT167dj+uy8iwHN4ggWGSE6hskMT6/Vi8xaQvBsBB6YFuA7ErXO4GsX3ty
y8cR9O7ipzySbCiJQHCttRhQhCakytnwrrvh1bJEbANUH55DE8UvCNB5BzxraGbR73rHVlMiQVEV
WijJluAYFhpYDU7ouTxgQec4b7uTHFfKLSIdzvAhDE7dtMessCNzCGM/2o48QcAaanaZtoAeg5MV
5TGKIXYjhjjY3HRsUvUD9LhAZkaT0Wx71KzZ3I4A3lmpUdsla2UDsN39nwLlVXqJ/mAmDrbuGMSf
kArOaSFZ4WLayXHhxiDpnz8GUnNAAN6t5QkXaR4Jn91gRRSzUVQ20SeojO4MeHzO1Hd+87AYfLXl
7k38vl/Q2KHEWHQp+IqWvAi4whRdq5BEFGB667W+NLdtBvD7F7dGaJg/LYd4jhooaCgFO3yYf2lV
3ZcZ8P1ZuoYK4xn8pRjYb5wQREMk+S7knQTRzJ/pycXzxPZfNikSNfc96FIILt4MQEbh6zSLKedp
BQqlz6/HfLy/hbqJQgwit3bvftuoH+/756USkY+Ehp+eyIBvmre4U9KtXLfr30J6wJXj74aIwOlU
bJGmaMlR+r4aqho10jXSDB8M8zEzYc4RtwlNjK22mhVfBeWxKvX3K+BbMI8r8/wWSzX6A4FvQLuV
XSUqd5n4C8ptiB2UCASQwsthHmOJszHG6FN2b62SjuTYSiU3hc7wfN5KiVSGZfsUTIhQ6I4X0Dtz
XMPj57OcC8skbuImFNCdQQk0+pVXu764Kp88tAiR1NYbeU2r1+TkYJg2q8PFv2IT8MYn8WkYxLpr
afu6+/jsxZ0F1kNy5pn9+iU9WaaQXhjhoOvpBOwUqFCxViIwWtfG/lIDUTPcdKgfwYiFMCbbbYc8
ClRv7ssghhoPyiyJ03t3dFA3EpOckrICH5bT7i5GNqaoNDhsvtXxcP9KyUaR40Sx1BsVSEWN40/G
Jk6Foi9i498HwgeMP75rpfln0jP7ZEXp9A7fX8WSt+hEHZ02YJGxhDwqG+uL4xlqifw5QZ69smty
xqFZhSrlmExTv6QeOz/vjqLWq428Spk8s2Gj6UcVPBWDtmjtJs2SZoS7MTLqaX+6HjOI69wp8PG0
vTNpsJTP3dOL4Bf84kELrQwiG/3SsFuA0/snlDiwpykf7BcdJfnffvPLHaPDJ/6IO0o9IpM9aaxX
CJpEovsLRNkGqtNrmoqb3KwOHZT1wwOOYwCRRAe/mg+o/S7qJEF+8vPgMoVRFQFDbwXttY2hlBHy
spiG80/M4NE5Cl3brDNMqYvUSZFdJw+h3bcZHFNWP+FJA4cfDC+vck1Q67YfwYy1DkK+BdROJvXe
0pbEFJ+V44fkg6liukWoJluedpri2gvuLyuVUJmws7Q9c0YXfKPjqrq1+IJBSNgWCpFhycPsY7Ue
rBvL19NwgFpioWg5S4Wj25n+m8MmC6F1AGNaMjo+FyrOCguSR2G1/dJd4zkz9RpTP+GAsfAssA6c
8IhuTKSJKpX9yxNMskl3u4Y16esghwgxYOPi2rnujv38XWsNOIekfQeu5oIdhyXqGtBtUwGN4FRp
yBf33bszGhyaKochhzi6fQg00D4CWD3khb59ZLXgGsRiK0vmh1mBboCuQKop0jgJ4m1hKhutwqBC
CU6kSClb+WNeWTYRPl8uTQDjMcBnU9pdnOf7ZYQ7ODGRAtWQiKQ+Ay1Do5xVIKd4epbNakVdyBl7
s09CxOg+Jb22kgBsSus0ooHq0fmHgSiEIHns0rmoISaB+YH1i3RES21TxBB9ScoAaGulTfR9cvMs
fqIv2NiN7heE6HPAkR+sTqUL5TV/dDDJwJ4C0CuBUcxMNQ039WpC0olZA/PPeYCaFm2fxQO4z0Oq
qCa/Bgds3YsShfAD84GQ9Qxa8p2iqsDCe34qlT2rmFDi0F+e5SaqJxEVPctgbedVAFyFIgsQGKha
1XRJzAUS8vBHrTPu9uLEsNCwhtj4ktWhSX0KpFunNcj1lwA+/Y4MuvLLIhDj75elXrIWV4FMwflD
LYB5TXx8oOTL5ITD3XJ0yDF+JpUel6QD/041dhjkOfcPvbHELpg3Cgvn7eQUdvsR69N1V6RY/b5F
aHaJrk7RUIyZj3BBuHITNKzQL4F50r3IIkrjchqLVUYOV+1AqAqgiIyKGTKThIM0C9RAG/Fo6lUW
iYZB5jF7EPcrqxj7PQe+MpuPgBiXxvEP10lfo9wtZ/1O7HoJ2BD4H4O2Yg6bBSHsYoFfFM4nLRoK
bxJOXOHvf/qPS53JAtxnaP0gxNH4BBlL6fhKmz6BwRqLGcDlPvCHOtnB6EQOTbj7AbEyz7An+ACb
VFlaKDXdcecG8eeoqJV1trrUYFoeodH3SsXdI84Tx63H+rxV0vyjdxzSima7pPeejk35KvtKYU7i
e4cUhk4nulfrVG5lsrK7AGekZM1RtmIg4tqKot139a4/4f5uXrYMxd5HpNWub3nTmLPJ4m5P2epx
1whDyFg5Ts+dnHCQC0UCqJ5xuh39a0QqiN5N59efNkZny0vWAJNDuHt7o5QptfNoqzFoGZmgTC4z
cDVUy0UfRuUzCKAMeP63KbQDETL26G17KF2UUANidR7zZNcUG8JQQspl2yfaHJ15/bv8LtncpgWA
Hc2+YMoZvCeCPCwXvBd1dKcLFmGpmKEFahvJDnS3Yz5lGpLKqTmm1LQJZtl/PuFCMzFo7t9QrsI5
JdKjoLPblaU/38mTR2lPQ83Lrsc7JS4dBX2vkRPWvJqjGwTXcpOAtis0eshXGApIIPYejak4Gs/e
8e47G6gxxZN/5EGxiuU83TfBVa6Q62rPcigsTRITV4x0YreshS+sNMxOsYfQ5pf4216X7SQBjMFN
d3g4ZLNNowTLYidc9qNlMneXVQKSVzLScXCNivSU0W32DoqWmPCV1tHQgqLWdkxY8nxIa90HJyp2
YleMsIZo8Tv2ABXp/hyY04wU33NSJrL9om4Zi5MGrJ71nGpYfgQg3f1HquiFDaxWJRrLMwjrJvlu
+wnIEAif7jMLH6IfGaojFmvmeqFX7CDldRzeNTyiQkkk3JmnQiyzL1oAi0cS4fAM+5/U5sqKcAl1
qfa3yG/2haWGV9K/Xf478+J7OvumYeb5Z2Wq3PJkK4hRuJr+6q77nBnJgFoxXPMAazzakKH88fX6
f8tGY0TiQNPb3lvKFhUY9+H0VzMLrOcklZNST2gmNuznm2NwCT3zrqJA/q4ytgwjC2N1WBSuaC9m
qWO4DkJv1tnFBEpyqn7KOdiBDNozYEwCDj6xCCIksGPwMF6Sw7pdAlmMAv2uMXtDD00Fxj8F4+vZ
kw4w89v9OIwcFFdhY9qOWKVnyYo8Nf6HqYybxkvwfrjYcNgHfjDhHSb6XQoTrwA6FGPr1AAKc/pG
t1Juvg8jQiJJ6r1SR44Ca9C6GGm3p412DEsd6JFNvCmZTN0b6Zj3pCpCZi35RLS4yRmouWvbiSK2
XiDt6smNvQwe4yT2NlJZRFOIl3tw2RJbVh7t57/eTu4bRRx5CB2R2+XwE6EPhNKmUBV4J2NdDy7W
GVp3SwVZTzInBYvLJDrxrpB3NusAukSNwZlC0AJKiL9pAmlwY2BhChUl5CaRSguHoIktPl+WsWV0
sXy0iOyBe1XQvm4oQV9A68cMPo/rV/a/+xGFIOqhC+xTPk9rb25mKCg+geMB+GyYONZTpjW/Es00
hJQ/eWgssFnNiIQ03OWimZvYejMVEeaBP0WjRDwFbzIl5YVucufcAbzPCy42gpyaRtMsmDCN/Aot
Wx73yJxljKbiwI2H3crM41laAXUuxawkHA63LCqft7uhdd32jWkIbYcptl0t17JNt2keWwaYe8ms
xc01wzmIHfFTKwDrfW93FvdWY6KRvcyPiQHFcfbJRatM7Y7LJaDf84gPDH6adCdqOlSJpH6FP1ua
LHQG/AU+UuNXKiH/EOcnkn5mFnJFhhAt0c+9PN8pRWJWBuLISNmft9sOdJuHVnpSMkd4tCsFEzdA
6POjRBHas5GyyaKK8anFZ5rqhpyDMBQYWgCMtoRVglpKg4YV22Gc/WdI+PZpWnUG6fQ8Pyh510yX
Zrc0ajKOeQQyniFM7jGacax/0mOjiycy53OmV249qIG1ku1NcY/7W2i9YIUqAEL0of4ftfEKN9bm
HS7mslytC3VDSRMRvBaSXMshiO5ORB8QjfqKSlolLcRLUVAM14iX8U4D5CE7ONGVrDI5sRyq7BVQ
oPEiREcDQVXZzNOBt0Gio2Ng0nB/8vMhosrcxZVsH4nqSeDbsvqZX+AKPKlA3ywMzIUUwM0rtkx0
+exXiQ3z8jJTH7iob/9Mn35qP+j36u6sTKs4jfXPhoNXkZSet2N6Y8qYPFRd+m75nGCV55c5XUl7
bjOc1t09i3hMrYLROJe2erdHyhI0jcLnySefbhwvXIIGcx/3tDHECV3SK+mdTZQ0rFwVhNJzvnQE
AWSV0RBDF3ZkGbiO907gsz44L98I8aZaKL2AnD0+4hlndShCMVk76gUsxjtDNIhfO43LEy3KkMSL
8atf63ALcmsloX3E1BAygNjAqCVPUb6RZS+DBaI4zb1SmSrVykNSygPReSY8b+AwHscC5F03OMlG
CZaT1vfxP4zaSZ/TbQAdGDgdCXmkj2ba/LV+h7q8sieKJ/dGLbofDCIW/ZWrpzRSpYq4206UlwI8
tMjr7RTjElIPPeLbF9Z3O7aEZjySSQnnWtKEAeieYVCRMrppDFH4hkz7BwOz3l/+3mfovPMNuNdv
LX7calChyFMLSwuaEKq7KuH2MYTuzMDx22/QcD0xS0pnOkSRR7TODYQmkaxY0jC2UzhuwY4T62Hb
uZlNtNh7RHJaoK+fXYxCRAG1xK8g9di2F2KM/ZYnKxtIWLdn8Dx8BE9LJ3V9OOtuCIQC+80+d4Lo
/ZEN2GntESft74W0vD426Je26fY7QYc0OkEjXg0yn09JGD6lc7ta3LhZ4nIXDAKGjj8GDLhjBh0z
cTkkeomyMx5+rTLOaiBUlcUgjimtuWUlrkC2HrDME7PJyOgTBj3lBiKfOfMCzE2rsxokbgkxO+j6
4u6HjBLdxg+83vNW5bHCxkMspAJ4bi743SS0oOe6rMoPgGPcZmM7IOzcHjB0g6hxsAek0ZaOi5+r
5Y/08PnMwWhEPR4qNS3wOH9ABDd98NsuaLaMdXpHEBK6r6KBNe6ZVhhcr2tZg89OkYbf1IkKpNgD
9DmJGZHoI9OC9mTOfbrhs/cYnBXxAlGV3llQsX1wd7Y2ABRPMdKkQmShR3oDeeo+jA0G5y3dpdTL
bJ6/R1hKZbta42yieJfZBFK485SRjVZoFjkJ7bIy3H6jInyMZXWtkWCO5ZN04aevwaxkJRuWlkCT
KiO5O374RJWpQ8407LwbgZ5+NKxzNnGUhZmWlvZ02rv/RBAcyaWOX0SY2PXOz2VIxEFfCUNdlXmw
PHXbNAhe0TTrV7iJ8EPqmgvm/YZDrNcqaTEq30cApm7UJxc9LgdrZHpxH8Fhx2+10F8djim7mmvx
9Ah81/gGfzmUpuZCEFm8ZvVLWD7K8IVh29q0eZcq0Ng6fFpyyAtRS0fRSVgjzuq6Id1SRIELO1io
zVneFMdMNw804/g+5IsoL2aOlO+YhkkjsfmRd2luUo8OVsvZbCqpdxvYqYmr9MTL3gdU1St9Zmwp
iJwiNicqTLmcBeqHYpcxkdmqguyEF4JLOOGcOP3S9gIvbyZ8JA1k2bhwhtaOqgoXX1rAU0Hi9W12
SUrBuVvAafCokpoqW516FS07z7Z/s1RbfQm7/ykAwxtCh74KbZwwkZMPXEDzzOdSyovxps7fsgVc
p0x8J/z13U226mut3jG5E06OrVhty6fSQeHiCHrV/4YFtY1TDB0RyPprpYtDkqHiRCVZp6i6wxO9
Kjyc1obFKrj4qjezRrZjubY6hRXG+GmTNUBiuhFD79KIa5uM8FUu/B0lmM0//MLAtjEKoQlDFIMc
E6hdZoFTPpV5KVK7Zuk+SVqrFeOU/Pur3uYsbIGqkogbuSlGZNBb6SpXvGmgo8hjdOtF31k5/JWe
9JjqxdtMMNx0NouHiXUk8MkxHx1y9grCY+iQYz8Ilwj3CohGV2CnJGtHBln8p4ARKYNtJuI8xTxG
oTckHfNnaZzPEAqajz1/Oijq3E2FhJcMpjLLXg2GrsaeI9x+J1M1uqPVAtk8AtoiMJy6I4RSlfE0
WZ+71w2VuQp4nEuFb7WoKFhpb+L38uBreeIB2DMGOBElJjx2tlLFh3wpEUEpwDmK/dvJsRlbfrEr
qInzfGhCGe4ED9oHFslbkpU/qmB7vUgioqYb97NOZFl0v7EQV8FhpjZhtBlTstFxfJKQhexhVE9v
MLz/r7RNX1AQJQMgwQw9oT+cmkflV+g9XgEG5b9lmH+yrg/6DVZq44DQ1rwpbLBjrvzGKu23Zfml
gL/Mrf7XO5Ba+gOyCfAiYRxubvWMYy3cmpJHDkM+8WjZbyevpTsa/qoKU6a8OaBV9KTSDapab/Qu
6zmUZpFH+lSosDp31jmTomkymfrhiCMswpK6pc1O3koRR5p+1Lhq+g4a6B15vdFzcyKGU+H4UaVo
G068lrEnFVI2+hKJD+6nb3EnmIRz6EoYGzv5qaXvFqcEjwEdwYXg03RpXlDjJD4CuJxpRGvJWyap
Iq9S5Uyg/L9o9Bmq3RWK1MlUGcuI+rBclrRwDDOctdl+MN05YH4hcAyJnDVVh/Lerl7utoqOUeyz
0LCGm9uItzvE5Wjb7CIHQILdfEDMfQD0G/N1dZhGcz7pjNS60ggnwmvWx1T6VCruph6WE+QYKh86
+e4KLpeIeTPaK/5LfHE5xEHlKEUbm8TrIYFy+RgzkJAniNgOTcE6DjXezf8O1qiGgeFtvBUzsG4p
waR2nY1XuqLyPjIpFgHeXHyrG7KpvjAMvLqkG001KnvCkXEhQgKuqmJhcMGu8ZJNEYn0y/5aOqLz
qd+0tvEWAEuqRPZsIdIwwtrxo1rqQVB9XIiBbm3PIWVZD756ZYQ+181ruI3UC49NUo+OFTV5VOo4
UjKBqx4RdXWrG7bG36j20bCXjQMIasiAmkvQ3FEJG8hwoJIwMibEli529Erb7XoP+0qb5s7H8VeZ
Odgi3qd8PBz5iMLhNBnAwIMnBFhc4uFFdK0Crqo4CAzggSd/gqPIayidfwCc4tkZhTqU5+UyGlCz
4sLVQO1tlOVDomLo8BSpGL9vAIY03tVUwk+qiShR1vFUzYUIJ5gXerfTmaC/WQicEdPcy9+WA8jQ
pUTNmd0HL9AveRAxAKG3o5ImJHaeDGAQyZdku2crlAg3Kvaf6jZ7XNUgodCDMfdYmlj+qltPR8oX
3LTlNCV6gr5/ZKKGaTCqgyJr+638ffhReBvja00aPLeJnYwNWOUsU7iO5CR+K8Rmj+1hk0dXf/my
OHUymC9fDKAEKPGCs6PmT5CJx6TvjYz8fbHgqpRj4ed7IeoHGVfJFcMoi9Rx4s/NG4lh7jK3ifer
kOxyfoRcdTIndIwbLS5GfFhpXEixfDZrvB7G8ZoscoQFo3yO5TfN7TZwSJW4PICzAkADmNGiKvhG
GCHXrrg8URCak9L1qVAJsK3SC2/2jhb647DR6aJnHArN3X0ytg9lDLZ4GOVmLQonXEjNI1y6w7h9
kWlgxSj0al01dEYBareQGMRoST5MFs67aMH0RIQGJowiqyJjyTockFsMsTGsecXmyWGFzrbjGqii
Nw8ktB2F/dcCKaAvgZalR8hOF+WHAbWjMLGhdglilGy2cV7L7GAAAF8JXhSIAXn51Z6VHyA++T/t
Z2A67gYWsl+GY0e8L5qI9fNDaaoXViZpmvPJZxpt12IqJijblTac4aADIGf2g5AkWV0O0PlQeESy
YhkQ4uskAlqQOPQz/PKpt93TJ7m9g8fhRxNoq+gNSJhv98uI2C3MA93s3oD1YSxuUNYrXfrt84I+
pOtdo4JwhfrkNnMVkD2VZ3PPGibXUL/63wUb9tqatul95zWKfFHCatHBR961ZPm0Bb+WhXsgdHTh
6qrNGrhI1yxINRraqRq0MkNnpiAgBW4cGyPg073V9SpT0qngqX2X/8/hX6/RzCACyz36vKsCvDRN
iU5IotGmY/h+VTva4D3rlFoz/ebst0dX7svAzHXeEvmi6y643NJa7N8npkDRKQQbkTqeRoyhHAmH
bduW19btGfGIq2i3VnwA5rXL2bQSuammqWRbS4bcmxrsZQJ4AjnqiL3gmQFrE/OVXsQlHmofzs4S
WFOJiNXxo5mLuztj7k3czxZhYNvoh+LEh3B3RZrZxkiTrOMLuQsbyB2aHG26Urq7QwDCe0mSBJhy
84vESLUTGujmJ5x0EPLS9w3VZTgl5HiDEBZkqzu67kWEUp2pXqXR3D9L0pnVB7dKsXLhrpXxEvRo
9DxEnBpUAD+ILU2MAmtiSH+0SLx9T5r4fXzyKgCDG+dYIpgzRVVZ9hXDrp+WV45kinZadC8twJWJ
sOlS2wWZMh8mQEcjmxZDLxY7TZzPul6pzicyj+qs+pDq6k1hEXlqLTedN2Y+kmfpKtK21D7KA1AJ
utrG7MFbfsjQB2xplMc82Z+uYIiph3qgU6IfBP8u3DF988ou0pctLp8IBgSMOgUvpO7bs/A5xMBw
7EJ6JF8uxSGj6kJgKJk2DSVfok9vxVDejP5c80GY3s39HhqBCRsyiP8oE8Uy/MiZyElBe+4ALO1X
hcPtudNTDSKyJu8s6hAdICaqCyl6vk9OJZPEMx6sTbOoDm6fcqpC6KJMkFO73MRLEEZEOTORR5ph
1q80wNBU58ySnsmN3B3/GbQndGga5BL9yByBkg4flb8dvkWX4jzpwsunKHrRQtTkOyPDstAluPKh
+zDeXtsvDW2m32Q4AA8DuOt4zwIIquFRof6ly1MNQAbPl7qot2N546B00ET40YDZHtXrTN/SahUf
WzZYNnsTaH18n6imY4x+MSYcSKlOStQNmkWd3rkouVWmU3tBudxlM1muOokhB4lVoRXwLSMWi6bk
fuz6Oh+jOthzwx+Za1SyFcxpRycX7Opg4A4pYPBOlwFah3uP5WqohHEYm9jYF++HDDAG7IfoJ7UB
fqnafnnnUxzZWUwrcMZKkA2R4RJr6I2Gu2/Mr8NzakFx+WOeiDBWjs/YGIDmR+0I3GkiqWVwlFu+
yUU7sRISMkrV3ARLS513vG/WkAClpDiTkiKAFJYCQegI86yAEdc7d3njP4xcq+KJq7e67Y4doEjL
O8fkjzTmS2XAB+NxiiKZ1Sr/UazP/LgZH15PJdVS/Hsd9ADtB84pvVf0SqGghYT6xF6rHw6VIxqH
nZUfUFT2xcvFDSOXDuaNtNpebs5oqmjPTUVwVE/n3kfL3ZjdxQnUuJvddzdYGw3XqW3EeLkHp+Ya
JN0kVjWcq2NcXnEBh5igHHymPgSHZ9YpkBO69HjJLLO9AXIVAFlmYBxVQKZtWlCZE7dyGRwAeVSj
G/+cT3IFO7lREti4FkrHRNmW724lY5vzrUTqHr9zyvFnDp7OY/OvV0mGlPEyiNZFOH45xPiCSnxs
rT14NiGBwU+wsFJ03mZ1OL150C6v11Tl7sobLXFkIUc2DPA61uJ+BvKW4T9AXdJjWZJ6ygEpvK6X
tdv2Dv8+9NWsqL37FmOn6DEkqYwqtwkubZ3fScRbZgPIMRLusP33PLxUsFLoEMQeN0nvjiCORVTR
T2ZhKByXCqlnDO7NYQ4LwC9ZgvMlgiCWf0Uh22eMBqiNco+RdYycS/XlmMe8VyyoPIyvDFc46I3e
Jpht2voddxaxcQOpUF24jE1d1vBGEF1WiF4kFWQfYOcS+SKzGv9aYNlgTfTtWZlGjNlGuFt2Epdl
JG+63zPSXSONAjO5EhNRcl6/4JUydxoyYJ8K/Nkr3BU2KGyBPIOulhkECiRhIWdcxTxyEH0Pvid+
SHIiBpQF6xAMR8slRLAcfxdf4+VOUTbdmFNp91z9Yq21yE9ejShTsO2zEHqOtXZUxDS8qa2jcbOo
ua5Q4GQBLvfh9KtjYyIFofig500e/iFnaSckhTqIx11TNar6oVvBRocCLBqCkI5IUuVzaus66Nj5
0zQx/qPK5F/YcmuwyMhncXWLw0EmgTTrYOZezZbf9070EhuGiodiweHrgsz+e8m8HOyQ0vT28BY9
ZOncP+oIhkkDBjSrJrVRor46vreins428i0N5UG9ROanpT4IALjgeuJWdO5ZwFWKw46ok/5GTnCe
dbQz5uw1qTYDAJgqnHx/QWA2NyFP08t9XzeeXEy4Hsub3HW7D2ttvIYCVdvFvaof40QLVU4MkUst
UPEpDUYTIe6DDqZbyXn5xmKdJ9D6bmbLfRiV+exe7sRuTkqOK+n5WDKItkOGEWNbR17qYQAnqwuA
hRUI7KrOgxMqSSHjHBBoOx0n+6qoanq+MUnztuBPNEiAVVQS12EQnF/4waJ8jBijME7cfF46Gcfq
ThkKBYatpu9PCB0wEMLNl3WgTSlMw3lRT8xQ2p1rDu+yKKIkkJ6ICcFuAy9SzbhlJnX/O6iv0m6U
41/NHwFFY4E5XMTj6jLP3RsUCbgwtOANTSdvjQFxIbtylQ9QAapIoVUhQxd5+lgWxN42lXfyWedk
b0xmHvG6zB3Q9TLvaZ1qcqi+1bSEvcGS/W1p0ogwrffXe6tfE9PDQ/yKi1bgbqn36ln4z/5K6dML
rYOcyLVpatjsa6Vf/qlPbIZa3poaBo72KS1Jgko9b5i9hWTYuHxJQoVi4ruY1Un1EkN75pHU4NlM
0ixoS6o79MCdi/cq0/rbiWoEMSDcM2q+nY484NrpYjNJfSDF6usqcUk62UbOz7ICFXTaq4gXPW0X
c7D3TcOSiOuzCXwTnJgqZIRshgo9NMGHlP9QRGvOd6oFZoZk0JExiRF2vHoLBP4/pRX/tFGzaLZD
eugZ3cqkrco339h63nIvxoHnhmVIP/FSq7netBxnTmrvi54GBgPA95B0ogyCc9zhqQg+of0Lv8FP
GtV+MHNILuOr0qaSjxcSqV4R1zcxmxhEhplD1rjt5RxnIMstcjGyZ3ZScfe5a9tfXGNyMeiPOfMX
wSsn8j0qpjzSwOcP/Cu/Wk0NgAFGZLUjCnEplrSvN/X+iNXIOAVLp3H5cLhjz5l0gKE81Q8xusQQ
0niQRgBu3toojj8CIkUZMV3wkYnkHRxjRb/prWY3q1oNNeRaFmT8i0Dy4ynN2/LS879MEJfLMEQf
rSfaX/eKSh4YgyhYRDSDonSowhl9zYFZeDVjefkEecC82NhjDGYkhP3UnQY2lwzJT57tleMiBiMS
xdCmaWHNYwPwwuWZjezle6LFUcI5cIqVO347VRETj6lrNdrL7vfnoSa2XJdnp2JF34CjRXeaBjoV
j3JfCRAm1kKi9pA6GUlNRPFB71hTLPnL+zfmuj87nOhN1o6brrK3gC0cliEW6ao83g/3Z4gJI65/
6XQPvklm5SXpnaXhjZHIrCVts3ZQbUInORks4kXBM3goI7w8NuAJT4bgttlCJMr4Bvyg9BAuZq/w
fnzAhyTYqIGq6H9VzJjYTvy48zWZyUu5QhVh5Z93FaDkafAgo3PTr2Z2YiKAZS0yJ7EaJgJf2XX1
gmuRHkd98wisSjI+mLuWBwU7rr5Ck5KNfdG52nmZgPogX3ONYQqqXWbsZAEasEMLp3PV7IpxG7Lz
zK2feg4CnOmzSp01+9D+O4IEH9zM+kQ9AuRs8jjAAcuyC2Hh5fj5+B6Wyynm5tR2iXv5b0rnKiVu
4MWB0dwBBEbQed7bOWYSsDb1axWMyK4bogBME55bd2Wq+2pQdds5Yvt1qYykle9aqJZOnWjDQap0
F+fbJHlgxlSb8dDt7NnXjufZEiW5uYgEfYXPjXrypt/MocNdT21gPNO9Yz3P44/IAUTy/8FDBhFi
KxxeDtPos9YZv5hmJD29jxRZvLNG2ZdQA8ZZ+8JKNWpMDKr7sCBX+a83oxne2mXS7CcVtaGJ5NOW
mE4mrRaJkNMH8WqM4+V4uqV30dTxcKwljlDUeVKUr7mvADVCG2YOu8d00Rq8wzZ0asK+gBX+48KT
YjQpZXKaLpcxJrJPUjOcE6SGDNZaidwRSedbEI0vLPAnBEhfzTZO3AFTkSOFXSSNSHY42MFrXY34
gUPT28NvMM2W+5JiKMvKBwFeEbEM3ufBunrVX7sS/217v6zvTEBb5T1skBvsEzPQaPvtB7e6zt4l
pK+JXBtXQm5uJjG7gqvO9kMH4YXDYUtS8Nxem1c305XlGRFtuTAasKt/NJIBtH3aLMVNqJ06AYg6
fFGMzIM0/nngdNoyMC9doa1OPDlMsmwZ3l4tRv0iB42p3kswabfPEBWdGq3hKrO/Sjt5OTgKHRx4
SUi5S9ZzlWtIuPQAsIXGCYCTArMkvjEvQauVqyzrKvYZzb7l4JckKhL9aVy+TXqj/cD/2Ax7Y+Up
lHrCFN1m+Jp4ftXXUUThrcKYKrIHqlviY8/owonSGsO1DQtUQqdnYl55zmLm+jVAdpQS7kYrTD3t
KgzabU5GsJqjrmUxJorIFLUdiOc0c8kfrI7SaS6+f7tdXIMQLlQUXGDxpXyyv8VVWSSig0e1H2+y
V8dm4DX6Z9gwv4Sj06wHj3N6DSqB1OH5w5d7X3l/8wmApF81EBqsqRFUFHjXflv9xIJCP6SoB1hs
RA3gWx3LlY3WRv8mxhkHUgJzkOGlCe6oaDBsFsyCdhUQvEkr7yP8hVYi3t5BPREB6qkJ7SwHqNSW
FOs9N0zB4zwzX5RQ60gDRsjz7QVKRiJyEgtHNmKpSjtvmDjGZerWip7np6u1EgJ5viqyv0rkX0cp
AeIDmw35Ww+VjkrH82yXMNkPrb3KeaCSw+BMLmzJoliufLeYuAs3VseQ+uE92OrJJTyqI06MZrlF
NBn24ybupTz0vM1eATvVOGff8P71ikkYAEIwnLK55RBekz0TDKp2h15rNAqRxwSlMIAAB8OCKNem
k75P8Z33AhRvrj4T/nudZXweGC7dcKe7JIv7vaqoHQNVp4Q91ceFe5flKQRiDGIrtR3ZkW0C0P6b
K01NlrDdseKy1jk5ACw7mcf4M2OwVZ3cHoJP95025nMaQd8so0JgaaoL0PIwj1yT4fKYMZBgoves
tkbqio6t3Bu2krMzLa4tmUNa2DutAgM8BedRUmtZ+//TJXJRewXAimZqE1G0+QpH+K9KfTbfb/1c
VWunyBiil4otVojlX85TYgNsx9JWTZrQzDGTm6lNGcK4TgXQQ6A9Yq3nfWXeBg8WL8dM4amXyZ6B
bIqDvsuFIEDrp63ngKi8oOxK7DBITbJtfhtkwAUYs69RsyfkbwdRx5tchk2tDVzrVdYWc3ilp540
Brwrz/59HjMCYdeXsvSBlk1HX8tcgYhk9QbXC3dZ/85RsC/8LUrD/yDE/SJRpL+sLTwn4qqlEpKQ
H2qtl16iTJY2NubxHabXyYvMj2SlWmkiG5IejNSe3uzB5FyDFH7KyuY66HUxd+WnlGX8ULXFM3wm
coCg59MFv07NsZAyH7//Uo536SiKg71RnD5JtnJKiq8val1L19uIp7LFTD+Zi+mQiSrtVOWJupVQ
Ak+ld2SvNIln0/pOt4yKDSPU/tGh/1vRM3XqEXBko+Dg
`pragma protect end_protected
