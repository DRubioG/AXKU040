`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
beXsS/2nG4CYsv9gFF1Ju7Q9dosqOYzztrYxhxxn0mXciB7k5CdesN1OJIqpJl/OCGX10tXIDXVw
+wPpyT153Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
APFOjVo1ZohPQq6zetOUea8clc6Me2xjHl4m9VtHaWfFdfZMVLK2sjR6Zd+XYDvjPfrT91mDlYc2
txPX1TyMZVtpfijgMWitfyqHpEzqcEAEl6tL7QJY1ivs8g1jYL/u7rE/TU5XYizUnbkNaR7ZJpqU
fl3tjt032+xKEupgFYs=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nfLqxBplOtHvzS30bZ1hKXWVrqduKE5Qz6kUnh4/90TN1O9nDgBouE5GgxkwHWhoczlww77uzAWu
Qn493TXQYsBEpR5BVN6Lsm0pTNJgdDP6x9UjfAhteUZuEhtAet0Gr0srKa6gU4FT7Q8HLwi0tGMl
hYqGiChovgtmp8VbRmEbXGjGf9LPLAdkVGbfgfKBj94b8iTf4SnEcS3K/ePlzxKgynii/u8QMQki
hxkK/JGORGyGYgZNNBKlDGutcxLfB3YR4XzqpSgzoX/YCjQqEvDzJ7rVom/AfRMNFT4prwtTx3+3
6VxVYVJqrAGWLV3CSvM+YbOlsuFsaSy+ROBRWQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Xx1imBIbBiMwpPm7CF0u8nZiZfvyzGo6etcthzPbtjTPeffzFoOczI1mx+eRGhdKwdWAxHZCaaOJ
0FWJfefy+QqUiLT9SKt5o4+xbxuBhs52X1DG/jzoa+yRRqPLRK3U/ICoHf4VYlNDgtgy7N1va/GD
kSGtE8oO9w18lz8b+TivopguHtRTopl5W0idNodqHrQwR0V4JcvelLobwH1ta7/ANQGPDTUhzthz
dJPV8Ygp+W86DSvKzS7EnnmsqkX6hQvq5Qu3ZRU+4haYhQ3cqErjnDsp/mVP/Q/vsDOmsUCEfBss
FL9iWxeWApkT8Wrfn8b66Twwx+gEFrgpdFbU4w==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bb9LILWgV4A8Tkng2uerPJhaRFrpnwESmKswLBZChKRHBBgXNhbsiTMp28mFBCVdJvAGu7zYX8p/
IXxhaQe1hektJPrw3/zi8/Kk3WTGSM92oQiCy/TqXbtlDfTk7DdZjNrIRbQKO4ILda5EQX+k5edA
GMFkzYTUS9hVhJeEQ4O1+uQR5DjdWOgK/42PlYGYS6rhjij6RKs2maQkqSoDalcg1X6y4KYQbxCI
JGo/2w/Rd5qJGGM9TXm9aMrJb5+dyCMXGsM+6Z1VbPyhbmc0ob/5F14GhFL/z4i3PExEWZrr5MLi
pNSHAeNSUFznHqtqjhTBPQCB/sFwF8rEylGEWg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VQlrbbJjaZTBF9eN0eEreX6XIsIfbuBuAnm18FzS8KhxoV6SHEfiGDPO9ObFClmNHHO/mrVlNhHZ
dr5TEkL9ook5rMD13SR4l2EpGzIcd3Y6PTETvGFQDAGYsk2GY5IPiPPbu+EpnnJYlY+3X84PxILJ
5dWX0zyqOPNWxwqqwx4=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
M+FosAnGvDtntYB2lu9psad2sQEqHiefEpw2N+y6YncVW3Lxs5G+BZsq6xBqeA33NfA4bY327zYN
gQUh7iKx4DjxkI/LJc8fQEx3AbVzbVCKeI7RLzP6SPNucAJ3cUjdTpCenpgpQ3iP7EU/zKZrmw9F
hTVSOWMrW0ZAHtW0nKwrZPK1apBxx4LORCnx9e0eOR70qIohg9LeSPZwpZF6pHPaX1olnqkjX5Qi
Re3wloUG8VnQWS/3/3GgwoXkWm+pSSozDWr9+56t3sBWO7YXkPxroJcvJG+jn5MoaoUZctu/fHPa
iKROh9QlFip37f0U8XKnlwGP4QBoDkXzQKNZMA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
5w18o2OTP4I6OlxjbXEJXCaGxtGQw9MzLvTtAP39EfTGkk7CAAJqVuqcAvUwgVIoTD3yYQ1Z145D
slLuaISr/frTM2/msDR4y7S7ssvGpF02UldZ94HXG6X6L7VYBLi46JFDPWZWPDh3KhiUMzPe3JAj
AY+BKR/AAxafmJzEp2yYLsIU4w9MZbB+vndKIRPgbIvfyxOi+xHCMr6500AYCPWztaUzXE1tHEvE
fKPMx8s11OrVW0zln/QEwDUnm3okLdkEyaD6SnXdwnrqZkXk6Ub9UbiURRWnP+0XJ29CoaqC0VRM
p8ubWYiCWdz7jqdB8psEX0h+NoSjWXH9Fi2Z/SqxcdwNYDCi/S6V8NILApMttDyfgbL/y6nt7tgK
DXPJSOKP29wuoYpwJ7bhJlTptlxEzb18J7GGwioed02HzVYuJxnhx4iQ6PMpVhp8begR1EA9lKkv
LzMoykH9W7Fcu0zlB6Ihs7SXcuQSnwxkZ0B39BYgg/El5GrqfZ5xNbsahlZyEzIVvlgrf5/wRJP0
muKJrwdunixid77ZLyoQuiY+glt7mTiWtExcAUKA9AqeDFOwAPRDhRIco5i6hzs38VP0JDeNXGVn
Ag2YRyiarTUP7Fqy3T3UJjObUzAZJIOo8L50Bi+WE63fxdVigiwkABnyOlI8FX8RBbGdxfHyDf85
LoUOmklL4tjMDeh9ZnTd1ha5PtcvGEDcpPHQPEH5SDlsCVn7qFf9nKs8xVRZbau7cwe08xQUQQPR
SO8DuxOSE7hvTnI6ovWC/EoK/095eZBSCkrkHTxmvSh8ZtMR+6pPtUXbv2WtkUxCo6SPtdUKlTYz
6I0QdEN4TSZBdgAHt0kjgvyUUQHFjBkL6LzLq4puJYXZF3gyU5pXemof77bS4z06PjjWVIdgoUS7
2drfvnVa/oSWFXHo/yOemcfdhTlpBfkplyn6YGJ+FA5iKtd8JW4f3J6JoW9taulT0aXzdAb8kyeX
rZfUF7nObZZpxJGQj2g12sQpScH+pyhfJZ8dj0mpwobktMhqnB7L3G1M8vQawh1v7BrLFrPRPyzg
mALwQ4KAW7duXt/Y2N23Cz8+93W+NzDrlJaUJXeVW376Qin4mh0H+j5Zc3zyuHJ3OQnhjd0Losx8
TItV285QBNF6emPkmwrmRQuhGdoFLBN0obINb/qa6gcOKysDrNudi5OrBYhkxMWWWN+XVvEKeb8R
exHcekvRlpGWpnUUiaqyrB9CzkX4M+45j2P/746Vo99iDz+13idKmCD3mG8DL1zLGcqHrLGFI+Ah
LQ0GYcD1DYM2aLoC6r7Cm+nDGdjUPUhu95usQ+RpD1CU8KFHmUklhyv8PHprxfhqsp2xMRMEgp1c
ifx3n5d24+hlfXM1vUnzxx3Zkh8IoC1DrkRO2vNrI2j02DnjGGYbdaEjfGKRKemp4LOj/C1DaKWX
uL+dwEC8DfQqKCdmfCvd2ewGHjk3Ul/hyv1enQr6s7QVG/GjzCzg/JbyaKff0YWq3oTH9nLhWrKX
yYIvf6tVN08P1joA/SlKgukWNjt0zpPCl3lycJmO79eU3dN7ifcq9T2wOwSnp5BSzluDWs7LJCrR
21e3kqOTbLdp4uJvtMLshx/7r2fbfp2ZvPdO9oaivTv2BZcEgAnH995i3KcUJfWeckr381nkVjMP
oPU7GaUUrZWZzrdl+e1qOh/0w2vzQgk569VjzRahd8bKNxxxTWutj795VsFuw+jxiYdN1kDVhWzQ
olZHD1MrBKxGvg7QBQZs2ovuDCfl0tY1hK3AvCOFw4xgeVCMWfEzi6vnDqru23RofuCMfJsxHQCH
MHF6OAs02/hU3V9/5Z0TvIDw3sAV93mpz2lBAIB/rGNs9Bz5rv1iNH9W7mkXe5UjAcsqJtwhH9Pz
12kU6Uv9Aue4bhga+xEiwoGfvmNHy9eDEDqgHazdvZ3hqmfx7QdX/5AGx0kgtZ6ZlljDSCp9XtW2
2PAYW+Od/ocy4BdUA/U+qOW53d4vLsmknuVYnBJ2UFWzPxOgbA237ud1m3DAyKuuWFki7kaiSZEY
1g9LwdsIE05A2K5YdbXm+mlNUZnS2GhBw2QaTDQ6M3sl2mS3hQHioAKxOLTUDf2xK8ah3DY/J0ES
SrFtwny9qAAZjoVlKgTp+tcpGG5p3aigovnGLW4eICnpcYm7c4oyCjx+wvuP0zfqcP7GBjgOseHx
d/6xfrB6TnLxet55AN4dLaMNULJ6Pz0S3SZX+jtXbjGSZ+IFXTQSzXaA+vEJCEiq3/KG0iA7pEY+
Dw7G6NnsKMzGxW1Q2cUvIvMqPfl9HqWVqeWhfO5oQhezSZ5i1agtcCjzYW8tuEyupjDoa135wlqC
6tQBAcURz8SCFoV1nJkbBY9P1Pb10zrNxtQPcFg7BWzsyA91XfLI//bcZ5vOqPN9Eur/0+qBc6aH
XDT4Nk8Jsz1BCjB3F2+ivn/1bbZ85FJZcj9wRxBpfdiVKLPCQ2DrYpTyPxxEMhz4eHhfaxJGsJL6
n3ZgdLm4TaN71Wl5A5qkqo1Qiaqme4y7W+BF6dmHmUD7epZdhTHb9juruBTccIjXU5zO79jV9p4V
rh7tN0QLWEZxjKwXtXWgO04Hz+YLqxzNJdo6YomQLxA5MkjOR9HSUh0oIV7LZXVzUPfD6rNhTJ48
T0js1nQVk9iQomeRaAWiRirv3R9ZheKc2Mvdz5O6JQVsvXf6wA/yYj7Xka/3lblZZy99AiYC3U3O
JGp8Ey58CVgBAZD6Arx478quL5xHZhMXNWAszKF9yXm/mpRYPj10ZPIbXSskECderPLiole29y2z
+Nm9fMhVTBeRhn1ujhKVrBViCighxpldHmOcigcU7I3G9bYOPP26htl/EHkyXxVQgDWjOoRvEvGf
FdN3PgT0F7EU/ExdRbmVdapYGpE22BQH1Yj74yvu5/vY8BHVzq6EXuQ4Hof0b3Q0OqArOUjZ7VZT
V+GbfgKeWMimbyGpMd6wcy9avJGP8pR0x1amwqrXnGP5QXLoBqPD4Br2Bjo5bigXElK3lV4+O6g6
WzL6gVGWnemTp89jrdFYGc27Pxmxb7zxA5zdDnwg3MpI3igohGfgv1gQ+RrsYpzBpAnKwZMmeOuw
lNB5hVsX9imwghlfA+fqPFACuZnO9dWUr/sGZmykpusYdTb4y1r8+CTCsykBrI/lnFC1kHM3uFA/
YUVMNLNAwaAmAdaMLPo23DP9XtxdFyZp67sLMQj6Se8kCQ84hgXskXLcM9Ok2D7tHXQPS1j7aHws
6L0ueHjsFs8dP++ebfuRj+UGHZ9movWWDLo5Ds7SAzDMMakrGyFl3g2P9Zm/ySYtQjJCLCQXHClN
z9FSKdXoWqsh8E3VwJbPvKu3Z6PjS+7iLG7zhn6DTQVXtdsrYAC7fMmBMwL3jIIdEhvbHW2eLLng
qP9qFlnGSGaZjsreTb9oovjb/dHE9xmZkaa01KP1QHIzoP7z8z27mtXWbWd6UIfCCcxxwQ9xmfKp
A/seDEAh/9yxcEY8ucC3IFBssDlLpFmAiNPr49+Vt7qUnd70eT3iqHq96k/H2WARMoSLEzq9fv+b
z0oHHQ+850YX7JmW6hb8zVXUKzlk9fUMXlkhg3DA/GGVNAj3S3VA8HHv8Hl9eCwjF0iyxiA2jsfe
TdATD822o+y9cS23hBn/xL1J9bOJQXoCMvJ1iofkVhO1l1LnLaWq8xy5f40Un34FMtjHSpdd3jWj
nPs7hYDDAMUj3RnEKj2KGIPoKGUHRdd5noGYrh7L2VOi04QTdrRwxmKzjD6xIxvIzehLo786IrIZ
4ECcm2i1CP4od38RAA2YIzzEpDz0qlshFswZRq6JUwwOUZl5siGvAN02JMCJ48S1C7+cjhT/Zz53
5ZuwJQvhLSdykeJIbYOvjAdqDfVmjwCmOLx4KuETc7de1kPcuLmgIeP/Z4TmX2iu584ZW5hW5/IA
YA5DqLCJSC1sOZrZBhSXk7iY96N/ZEL9Qgt1RrTN1SKhR6PtyaopvhWaGWq5AiBl0G2D+kLLzbeZ
i5NnCZ/MuqGR2XpXFkMKn2DWgJfTv3VoW6gpv8tnHhAgO8q9QxAKdtJrGJq1Ih5BQu2D78vivhbM
Z48rSBAZb03jDf62AYQaDN21gwZPdcOj0nZGY7m57hN81OrWRZgkYoKCBplpOjhP0oBL412j9Fk1
ng==
`pragma protect end_protected
