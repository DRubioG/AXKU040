`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
bCLM18CFa//LyZepYe7jTpZERapHD7ZXt6u3V6+KFJWGweIRYg9NeMvSX430Ldi8BeGy1Ba3uENw
bbsrWC2Rhw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KtPfdf++KcyFlKJ/x+05CfJr5wgaRud5uC0+mbVQYvsCxc9QehHNja3AkhGLko2tlGy5C8RLdToe
GQsI6VQb1a/jkLk+Mttca0FbvFJOpN/cbG3pHA7poJav1wv8BPEhyGGOm6vowHeO416XKsdQJ1sF
S5sBvjTr1yNDyv/bl38=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LLWDmTipALXnt4v9E2v67GiFFR+f0QcykPiFXI36ajYNrINol/aIJItjxFqexkf3Cz8nuoxpJJJD
jx7JWWMzTUzsonIsEA2sfyUNZuSGPNf+OPsaKL2Amy5KfYM2H3TD6uvH1KirZw9CiWfSzB/RTvMN
VL/zbP4EFfBXQ/mslsAWOK21KRlwq/n73tX2hduSHbBU3PmV9nm+1ESdyjG50lVZyQatkRW20Bgk
IGpeDAbSK/vqM2ZRn3pRkyPj7jW+KFrsrDR4eM6vHui0RCmAAq1TzyP5wnXEm0i50UTUySDsSLQB
qPzgx2MSgbfsfEIuyHA5nSo0zIXiV5XnwHJVqQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
s8R7Q9d1y1kFMyvg76QUC0tSYxA+vgtN0gehwfmfQbLJ6xJ43+vlmnLC7nEiLk7f9W6XiZtjoAcf
dbxQqQFaaNJr81moDjptTMGy8gq2ztJn+c8oNOVJFPtZGALxTcIB4cZiQZc+h2lOTyF/vXvzYOhs
iXlfFqDD+j87Rx8mnHq0PTIxJmK1anK5n0OMPvKwxqcQ4SWLfKV0uv6Zpr8iKsGWADMjkALZ+g9I
/t3HrpAaMYQKbhUzDSFZKILu+ci5IIQ905o1ws3tY1+T65gCVTQEte05fFFeHvk5EIc9IsYAfJKi
D/qlfkpxOeV+7lZmzEKq6H3o2aMjs/sgJjE6jQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
u8LNETGnleHCpa8r7CYqQP3oDb9PBqweo4KRh4Z+BSbklofkaIXsWDCWLubWse4tvljA2oDdyDDF
SH/n0XxyjfG9v1yQd+vpD5vPPEaqS0q5skUABw89e5ceGGB08uohfZ0col5aOJqqahELPxpQM0uI
R0nYeg/g9hz9BdzDEZuiY5MmMk+4d+6hr/a2CEtkmWBbfehyABVrQI10ox4UXb/YBfQ0oc7Cb/2c
+nbpiiZjGJWrfZ2rcNGhJmceCGfP33CozoCuRjAsW7s0RHD9ArKD3ilqMjC0Hw5YR62lGbJ6QHgl
cg1Bn5KN4LxtNV/vF3l9lIMG97FhhGOOgYBbCQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IsUjp8QZ5nLTDXY52g6GSAknHN8svOuyeqVld+2/exxV8ceWwIeojWzGxaHGCBkmVEbNV/LIXE3+
a9aSdx007y9g7te/Xm/xruWyQFGuJ/98Hv29KGB3UowweUlYtbtpYIBcgm04RiDqNJ5SFGEiDM0r
ltzAIEK05/pblIvpOKg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
PCuXJZ3+3ZGPxrh9pvQGG6TE6ZBpsBTSgb7ZzFotRKUv4GUYvZihoyFjUpODEwLhWtxuMtnE/wIk
3lix8iaxUyzxzUHYd1Hz0m9TYHeVDHAMCcKR3UxEosontkNHH9IvIV0BOe344wBANU+fCLi0IF3U
+e3Yb+ljFD17JLtQ6xqYcBK+oWQaEQk7YQUXViWGK04lYHxpbMbqI5i6mLJJK8NGSVIJjZVyTkdG
fAmL/Ta/BpFaBCCslBtsYYFXkPVsDWmMRVdEL3X8lm34xNRlb73OK7crvvA5CF1tflZtjeIj5cVL
ntO2rXg+YtxXcR92noUKFPtxVki8lq1ar9PteQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135936)
`pragma protect data_block
kQca5mOJvbH2jht4MbdVXiRLY4CTlsdi2guCrSE2UWxGQeWoh7+bbCBJRU7OVhjgOpr47gb/08Us
/fEUnHY8srN0TmOb9pL6tX6NDxP+hvcQwwKQ7F7PDrNkqJ6xz9NcghLXgAOrEBQ0kpy+/MjIJmv2
NDvvPsOsOez64RxujUUlC2vQ8m/6aO6GHCsocREPJCetwn/pJPPYi3k0i1uzbUn2AJKHJvZUYzC4
znMIioevqdhHnFFJkxhAP8Fw9tInrbGEVBai2DIfLh1fUZOLaKHuOp7OnZXcLkSuvfKGWrGRxLes
OWKJVl0nTfITNwfyvN86egvLrYj7948Nj8M9nM6/9NTuIxpSaaYfOF0yGu1hlUWD9zimyASdgw4l
2Wc30+6MdY2kJpvObFWka8DwIKa+0QKgyYL6rAyCugrFDVhLDSIe5aSV/xmabEmvsYaGMyM3C/a9
/kPb//9qo/1BvGZqnj+6kjdAYDAsnTYR4p4GRndwBFDowis49Xm/FixWSJSh//yhFVklbrDb6c0Q
Qi0IoXG14FImtB5JZoeuMlm6iZFwRjEEXZoN8LHuIX8eZOlcOO493s7/anhmx9siBua1KfUN22kP
gibRcjnJ/DmxLKH8Yh6YM/743FArkEFvxMhpsQiEZNOoOvgfSvpvNjNBXMlMY9WHaWgstzjVEjC0
GTYz6plUMqBpAmBgf+dGOkBKyNDev6vQ4OeoU9hnelDFrUXmhVg1l0E/dOo3z0+PG7ysT+6oBF9b
XZWRwRtQ3xJ090of5pBWvqTGYYlcuLvaQfJSAsPM5xvjqvug4BmdigOvi6VrO8yPnJRKvOTrK4mi
blTA1u11CRJxlQWH1gtS1nJhqrhrxzM200xyokR5C6NS4+3kkREHJEg0KsLCe/hgMZ/TCnfSGct8
05bX9ULyU/7uoJ6oRSDVeF8dXl5nY7tmCAJXo4e9k6WgRDMFKrbqZn1QBqBLsyNNm/KvX+MfRYYc
+x7/W3UYp9jju0LcCGoB3Q1I6mnDR5dnNtnS38Md9/RqUHr8cTNEtARabsgzEk0VEcFUIB53Nehn
qguIg7V+NQFM/Bw4p4kbwBAIKrTVN7nZ6oEujKsQWqI+k3zWmiQdrPFklcHWDYKphCx6Y4H/bRif
5OleykU8eXSgjKS0NmHZv9Kl9qPXrYkvdI+RKiROByHQpUlT0AenXHlBfXNLG0AQBJy19bPeRwep
jfs/GYFTAt0G48/B/k6oE8czw88algXl6kfdVIA7A3njQyiMHditVx6pw9Frr9PILOuhxAmEYZxB
Bc8H0ejeyj2IhDsJz+8bCAeGatuxoJSTkrOBF3hsZe4nIkEUJdf10VQP4Ud8N7AKIMw4aFNUNhPx
nzawoGDjMFI1lrVhEIdwJxk4NBs1D2nfCtR92NQaD4/cQpRamIT2ecSS3AjTmcgTjqmPd8M8P0Ar
7VbRUiGIhMj63dqxBJOEhsyMplnglUZPZUgsMbZpC+PZEj4FyUhSedxMgLxLP41NeMOChF3y8K8P
3OMu7NIogcvLSKnN1G06uvcpZah5Qinlrjzn1foChnu7DZnBma+nh7SciKWQ13+ozwKCLEIaBhoE
8qaoAaY8ZXsVKrDS4Pm2jxHi3GxmrQrsulHx1n6SF2jKJl3u/KXc5HRtwUN/NbVB9qsyn7dmNHUy
SeCYDpaMTLSShrvuhvato7p8GN62qwYpaRQb4wABuN5rTejYGT/aSPkvwfCKEfKtzwMtnFviKTVi
NhLOzSaBTkNnfZgCrk1Ad5tkufc/nKY1lHgESHO+TgyC18haFMgDOA4we7sabxzB3Mfgut2its/B
1Z56gupiEPDcfzQ/dXXswKESR7kVrlVGSgcKLPdCxtQfjOwxn5PSpnP1oByosjK8au8XCY69Cza5
lzb41NDkeNkSaWBux7cSXt9wHRfYJfSSh3qeawdMBujvARQhFIZkcha8OCb05zAZAWLBbVZIPSWz
WlMW3K2kbDPveXOq9NKnLdIjxO+KD7P4+xSXqgF6DdziAYzbPCxXlOgFi8WdlxsE27yD3fG1RsMM
DZzs7K4YGuFg1eZW49s8dJzhZmY5frbmD/xYzwzSHWKiu/MGtsxzDQitwPW3fWI9jGgCEcec74OH
mdFSqiUnYtdYcxoAVGvXxHwgsWUHOlTc7NfGLCQDJl8mVBKTsJSZx1dHcjw9oK9Wur3Qfzemq0gj
xBPBdYjpT9b445lnfQqKESKZ27i6uQilFXtP26Gp5dJZ+qsMm7taObCeWad7SEIimrGY4DsUxQ9q
YNGWOg3O5i/J1qXma3u4bgM5djDZkCjFWslmdu8k4flTol8e9XxB20u1LUeQ3/N9dIgPNXAHJ/Ob
olPwB3xiMkEy1AEJmHetvcQN/+slPyOdMQeFHDWeXYsKkg9BJIYwdAdRDmBnAGKoBvYjf+zDxH1i
E+Mniwz8BXA/+mRA9ylcXgxtI8GHuzPelf9fWCsuYC+q5fyfBjDU0HFGRwKhPz3sdU4dzoXCeD6G
p0pHEjm1Ef/oCCCvroAZZRomNNNl1MgDLPYrfioDdtFA+CJLsGVyd01uZgoab6zmd1pudDMAUcnd
SUdVHLB+Fg9P0UpcPT442sEB3rvGMPeV59PSEs2rL06Me6r9j/DmSEib56dhiAGYG+LvczphAHrc
Jny8QJRLb91GouxzMZpKhaPPdTfEPx6eG9aQP5Q5jmpBjb6eM7hB82Jpdo4R6W0pJAjyh5LV8Dgc
oEvl91bKF2Hp90NseD7YwZSE0fK49jJiQa7sVjKiHnf2Ict+oTIcLyBUXzISiIAKp9nXbFnAHA2U
11+gfpKiwivvHyTDDsbTmGvU/5oqIwgFcTzRNm8tI6ra8Ipg7z+wY5y/ARm5PE21y+TEJt1e8WQk
lZnDin7qOSKmoKPMihNrryRVmiETe9fRFQz9+sWbnuZIPo/p3l5XvfZdpYZT7E7spXgN/e/EiTZa
ZSMuZsGZAOfxSh5oFOyCJT9wvOKAr6ZWxSvI7reBqaTHDa4gzuO+WTaPUAYJSAmfmFDOc/GcD8lw
yBa9lvWY37/d62qcT+5JSSuk1qstzG1HquqzEtKtS2TLjtM/+Dl5g1tJxp3MB54QAzvggjDPZWoN
agig00kXPya01arkw3s2Mc17sx36i54N5em1cPD5OQr5XRygrWc+qfyDLaTwn8EVi6WaSi6D7pU7
/1/wt4l3J+19UlboYPPMotPTr0jtaJmv2SM7/Qtpt0srqUAnAzKgijWLSCJCmh2sdFqcx8PANpfN
inu7mf0wNlfmRqKo94MrXzGJY0qE319v0WnI0g7OAHmeKXs7g+aZO/nAuBJ6eZAonoxChQLhNetN
AGkG0QU7dO57wA8UfiHoQ3kQUW53qyzixxxBOJcFKMCMLYpVlOdsVwUtRr96T4NBgOdXpT13aEni
YWv+t5RyYHo6HnApo7KcHuU6zU/9JSb1I8TVV4Pr+FrcmxGLlrhThVBbDUl8VykBiPpznEE9/7gL
9rN7WtQ2VGoBLgbq1EfCfQYMFWi6ppwjyIwQMQSU7t7LOx5ABLwRmhoHIn2zvl6XP9IeYBP2bOLX
rl1tqqDqwhzKV5WjHwT2rjB3rfgTxnTaSTAldaYbJKeEpDAn3FbreKduJeUOKq5O6qO9RjPs8ZBS
5RbnjFhPbAEqsgYIBZFDKyngxwff/1b5VC6K0k8MAY3cBlvngtDNep65FaX8xdaroMtSOPcbnYAG
cibpXKV24hpe8PA7kOwNofKCXRn6CQoeVCa3bUw/UOf6xIbODHoGQ0+VM2W/GvrZQbnBCgm0ObMJ
TnAYYw53/XpOHlS3YIsyqUoiCn6i7RrzAaUFr0cT9bKliBbTzHhiKFl+JsPZ0+04Y0s42LMtmhkl
TlecE3O01RGHuRJXpelrtFBfSOAwNhWnmMjM446B+qeXbk4mlp367+IdVOdijqhcQ/9WXO4hQN/o
JU2S9lGPXvOws9eRja0Qmq7PHzED7AjmyE3dfs2t0g6jr8YO0qygsF58Ny58azzKUXTseCYjtg+t
alE3l5XgHrRAp4BzfHhKjvTDvChrhCJZzFQqvTVhek2huItUNhKVqNof+7PPgJTZfjItgvjlBF2n
HqbTS8U0fKwBnNm+6RTnvc/kRCGEV7AziZxJoC4BkAwjY4poPzm/fOnqWhVcd9Jy4ElxxEyG4Cy6
bmH/wMCrB3LIZxiwR3bE2J6crfv9g6c3t8WQM5KZttzdblKvwKwylkujRk5f2hqVr8xxFVtTpPdF
xCSb6CvFATEyclHE8y34AECeyfcxanHuRJ4+YC6jW+2AN7mw9CnX8Vj10SCOXWy2j7syeXvQS32w
FG4XYD/E8uURNfeM9YUvDA7SHFabmJMLhn6J3aWR//xkNSIZrqb4vn9BS4MhotOoQFYX8S3EAlpC
TxkD8qwBeUkuQeHLWAzky7TPILqGDIgMMeGNgv0AJscNWdg5DJWkdO0D1BHKUMh4Y4RJr8DxJih5
SSBwdZPVf1nW/6JjXWQmFLADrsNSn4faoJoUuC8m/ctbA61+Ot5sLN3424JsbW4imjrIpm9c/9Fk
GgeEoDVu+mIBnAb4LlrdQB8KKShZTZqgPoJKeL+kUgcs4RC/fRdAv8TnuKSq1yXaEi67N3UAF/TF
XrB1VGvyTMLTovvYbXZs7wnBT9LZkffeGkAM6eblhj8Yz3jB6xzAJ+Yz5qKt3xX01bMARsAoTA9X
qo14m1XJ2hvGfo2C3EBkYQGa3Xz0xZixGdFUE6fcMDyjs8U01WFq8knvbWKK3TJr1v9WK+0M8R1S
DSD2HEmjoPo7gzEkmpmNm6MhoMn3leso5irH1bjEPFUIYSFFXfObdK1DD9TiJXy2apnsSSmrz7Wu
im4DDGmF1XwbtFRr5SdCuJz0Oz8Tjcj7n6jl51TxNkn+XQLzHlxQYxknTMG7NRgmvF+Skcj/a28E
5wx5tmdlCjDF9QsiMUgMZUzFiMV8xZXzFD0jRGYbbVSchLYphtG9htD56NZ2cnMxlIi7Ia+N3Y1J
58eVpiUwlqtJ2jvqtEgIHOj17gJyxgWh5Q7TBOlHJzYWYLEAfw9qO/b+c1+hZ8xEua43/qs081MU
QFx5PsSQ9KsjmxezjfmNGJe0+T/ckalt0PvSYq6YQkmaVElNaA8hixwoo+MstFVRoLnDMKeICdMp
uG+A6CYZ6Hyng9rJZuBEbIa5/4KbiYebmIqt3+JPJvEh2uSiOG8b/cULPMyLYxUO3GtR9/ZrohXt
tnSeyOCwm/eErsB+3SK7bjOjwvkBuqXnVt26RTol1VwohqJtmvkrJ0xWKPDXd9MUrNWrSj9Kkn6E
ES0Y39PJf79GuqIih0nqO+BYBMi/v4wCvpNeflIpchMugGjsSUgqF8VtPT7Iq7aHvrCfjpcCH1mi
mCVXR+LUwPf4lOGIGhN3yAfh0oWcnZoIaifsouO3DXpucvXIWv39hSeoDzHS1ehKGWXvgxwcjvee
vG8g+opvEyuorwA1kGP5YwaD3Fy5sMTHu7nlZF2uGLYr8Gk9fFvTYku3h4byK465MS9RCsG3igcr
GXYBj1ZcbJiDggOu379GGWyX7wtUvV7qWFfI59rr785gQZJQC8PDUzuk4JXjSJj5XKcXFvKKH/M0
8s/ao74bHbxpYccz10zKth3L8TvO5W8c0vuxRcpEDyqIQP3XtkDNKGk2IZHdE5p52bQnLKYhPovn
p5lKk8nuj0f0AFAZOAvTn3Qi5vPzxPImF1zSrV6gei9uwFx0NzASUwSY5TWZst3rx9vwUWh6kxRd
XKP1lbN+wdct6+PhTRCK/eyJN/YixOfiGC7fd9t1Pi8AiSjjqvtFFnBP2fThm00jf0utfydN71nO
qKuDeveNdf3Zc4WoYch5fv3qnbGWRtE+9O/SsJX7X5eR9wugXlBbO86XnAaADMgQi0BLEl+eEUPb
4S+FMCRVkumEki/tkxZcLoaIyteS44eHnFogHw0ox+AWsOPqfHRwMBMk8AV++WZdIy07IewJoulu
4jCxvTm/GvuzLw5zioxJBJAX51/PxHVypBn3I+p7ImPWLgbVtNyzB1IL4ug29oRO/5ai5j9MisGz
bEPNAUiq39Yu1RXk6ufD6KJ9NjRr1AnVf60MzZBWXaro8CfYtY/gOC8BvyYrEBl48bczZvm5SN3p
5AHM5GqVM7UeE8Na4+P+0LsmqW6CiQV5s/yrrsh67AGsI5uRWhp9bJkdOzOZhgWw0cghIbFHCdqE
tb4EOIaUfDCEiHE0VopeKlF5wbyg//pAPD6n46tpl+HdC8q5IpPsk3JFH9QveM4rd9+yLJyMbK45
RzkaIRqQlaG0ieMvnFQfyoGkem5nmXv6FnVTMATrAIZRjDBaMghcMm5M6DKpshFsdmTAv/qSUX4K
BrYXF2pLnPRmwS3zj+mNMiRHs3Ue8l4l5g2RXk5Wyz1qKehQMa3X44jWJNSnNdFAS/oCcmYawo7L
an+s1KZCOpxy2rb1TbF3FCb/KPKQj6E8q/CyLroq9eVOEfBbb7AXzOxXmqdDeyCXYYIfw30FHV2E
cWbuzhrD6vKtfhIVG4yvlK9uPVAf4G3/uK9ODSQr4jA8Ob9XaNxGOy0Vh/XonzEi1zHD/Wf//i6g
7T+F+0odlOGZgvyKvTPp9+t8gpL4BW8WTfmpV9WdbLfV9F4NkRPT+/rmMKMasD9iqBVSRIqv+vr0
GVqw8LKG4IDUJFh6YsjHZ6wFuzJOKz2DNdAJz61rYD9poP6x9eRqpgji5JAbx2hSmT9DACMPiH+f
oTB609Ra4XXXgtEQ5ki4+8dXpZFFQ86oWRpjjz2IurSqKq67WufG8agydCGvA4nBri6t7fuAGET7
cPf5/y9UHC26HSsBISS2e8t4Cs6W/CLjVpTRvljNTnkmiriXgOT4+mDxXiH40giTkn3GWVkeU2HR
xyygnv143X3Cn3Hw4+puf1R7+3df5gshU7OSdOZUDz5fAkGRIx0oZoAMoPORZMwh8LZi5c3Jp+bp
fL8PJoMvKYYGJm74pBfrOVvGavE06zT8meBPFk8yrTYzygmPK+/lSbiy0cU0cEN+/eM+BBWci2Ze
Uo5p/OFIN9zfGEYXV7sC8xM04LDPACyMvgs7sfSWxttYKm4U61lzczMiYEMvEBo8UtPyMshJPSAe
RhLjIXmu/9WQP+jazmSGqk/40kPrbR6pkkn3er/qf4cZ0Kjzn6c1oVDLsoF6aTncKJ2MLWZZ2WpI
QPRHpW5Hrsq6DSFanuwZE6jiTEoNgovRZwaeCpKXZlT0CazygX3rNRf4wK7+1cm2Y8dARDwAcenN
ZJzdLhOJMLhnPTpYnWS4UxxAeGNxy8YfBdDZM3lGSh3eTEY9zkf+GsX3kg6T57v/8EsYyS7jVjTO
uSBBrOxP8JxoLyZGa1QFkjl8sTUrYl4/atHR7OjtwVfqlvp4IDm315w+jS6pA9bqt9uu7h+nMuxM
AkgdIpWX98Sznfr3EQCbs4zT2UVN5udAa+tzbp4K13gvg2/HyCz9cgmo+uq80HEFjVKNkk+V9eHS
/cezDhbDGtUqNB84Kw9hJMvXLeDdFIeM4Zb5I4WLPyBrny9xzAcpXPeUE7HY0Uwtl+d5L+32PkVU
NmMGYSzJehjM20Ev3MyD8X4wLBS19wpXMDkpeX9As/29lwqz0oMGJhMQNtYNZ9BjUwLpiUVZXPpN
sYZXgAdUE9vGyLrNOmvH2n5jUbJw/88UtXvZZq9Ns++iB8fP1LTXcmHhrAHb0Qcy+Wx0+9wD0d5A
eHqTits8n4xM5qHxqy7qD+r0KbjrLOs6ceNI6/27fZ1Z6Q8aJk2TjmMxKGui8qarg3RqQh7wD2M+
ZiK+f7Ozmy09AzroezgmwVnnW83MS3kbxmjJlNMz92DnSKcBeqIADuuu3/yjoBscZQfMkSKCBcBo
6PEjoULmA8vUXBxbjTb5DFqTBd1ovBacjXc+CJL+c7uxOOmjg/99GgdX+iLNxu97RDt5Q4cLvnww
Fwr0daM92csOfuBjcKCmHiEQ4lYnbkhh631w/FvEkU7tLz9WGEnANXq6lNcq2zmZvvwhh2yKWYll
IX7H4mUdS2rrjQzaNVB7IrXSUwb6MnSkLZS2cKpozEdk1MX3loO+BqC9Jbae34kEhNWWq488702P
XxFFa/ah6dhvPGISTQGwRkUDWHi3f7pSxfcoV33PfbpIHNwf6lC59r56RxKCvMtYanm10m+9PCh/
wtQCaB+K2XP1JbAm5CmZfSUPNRzkFhSUWTV08zrSw2fCuTCfEmshGyRD+kNypkJy2Vp8ughUrMbl
Iy5BR/irwkhOfQB6GZ+GUZTB3f/wce/635O77JOEPo1jfH6bTetkA7Kofsgd6fvGwpY0AXJkqc80
LNA3zelVvkQAFyIkuidGChvr4nlpvDHUKOp+tm9Ddy2cg6/kj/WDNpqCLhSx4+dnApDhYN6DlsZc
vSBTGBRamkoPJDvK2n1k4tW7Nz782wJMOHet5U9EmoaB1nfnoO+3ITU+M6YNBGLVrESPHpnKMsbC
iNhMj64UvqOG8sd2i8Uv+7D6q7ZpDG9DoLDeyBzNCg9OaSkmFFupEHD996zifyRNpJIQNPk1Edo0
yhu9V1JvOZd9rwjeKgGwEm7/bFOLi7QyQp3Tc9SO8acQozwb8Q/9vCJImUvaVreIGUDxMliA7XGJ
JwtlLcGqxRUfKbva1tRGUEA85R4X8yn2KZNmR8pnJFHetQUGrglGxiEGFglI9fz691yfkDopPYCG
FIkqwjoYK5Nltne1PydCZOJ5ZnqDUMACDfBCaUkRfK7yqqsPhmBzKfcINj4PH+8furhIbcz6dtqD
EgshgrGFwlm/Cr9eNcez9rMLs9EO9ZnQG0BoOa3qi/EnQ8JwQ/pUMNUWNn3lI6h+BLGuysKifBID
wlGU5EsBcbWaZ1qp5E4AEqg6LkwKYQ2bc0QfTloHXigyj/u1+rnOLWJPoOr9N8lh7OIy3Kt39ct+
MCbXLmAosTKEJnZPEinfuyJWEX0zmPUoPku+0niD1uBuLkDIXxEpBdeQBUCGF4TrXMo6MAGyUMfI
lNc/bH7VSQ+HdilOUrqnD7yLKsiiH1O3612vgTqP/vn6ZkhEEpXeJC7n5zbLV1UPxafglQWHR2CZ
Oib2lMfnxos1GcQ2L7hWX6vMMUgXWy9lpl56wXa9SrEGcoI2StrTfw8qyCdiCLV/x6Zynt57TpnR
NSo9Q5YyZqO1nobk955lIiVggMBSyd0W43H/Mz/AuNU/ujlflkKJgU7jpiAmJY+N47KzQy6aoDoc
DYKld5YuC0EjbFwQBj+izkrp2rMwZHgcV36AO/d801u3aGtC5q5aO8P4/G+1U3fLMzsDTcb34+Pc
KS3/6oiLjvkf6z6Z2q7oVi1QUbI8uLyo06ftz8XNXgRjfxdSse6t3rCinoKqTFaVMnwPg321O0S+
wTsVr0/3/fstBh3Avs3Jwuya9WaHnwMzgrjdHBxEy3eaEDRYYf66uZyNN6A8qfkkLNfRcsM+0QU0
ocaQ20/F+eFAujxyZxkdRkCYkcjhxKiPH/LA28eZf1LRsUaSMpBTZkTP9Q4B5MaNgZNQj73HlftR
0jqgQkXJd7f+yoKGD7xubSs26uhkZwSrhtEMzSPez/TWIWBz5sSl4rQjHLidaRGLzat3ESw7MDtT
K99y63NW+FMRLtPVIzdj9PwT06+1UMVlfpXXApDxfgYALjPDTPAG6t9a7benNAt0KgwPUtMbavzd
1eeqxcy4XVuzWBeA8JBglMSKBcUdo6Ks+YSZaLJi7IQaE6vpdt+7gAfsSLzfV1mOivFtijfjEp/h
Pj9rwiNsLq/R6nUBSS3WIjsPurZhgwqkOzax4unwMerHI7QPnN3J30/ERI06T/8vma1XlpqPxhc6
NoYuVglxJ7M7swrM8W8uBFb8sUDTjI95NSMATVRZ4KOULjgwcivUQRcKM1/csphacqpQY3P/6V9L
l/i8OzHr9bJJfsXCLhno295WZa1FkVhpx36DQvfKBoO7dUGwmJIBMxCnstoNVdYT1w1XZPkS63MV
VZgKk+ynUOdCVnf+Y9iScEsvoZ4gV0zQKHzoXo0rx1LDlSYuIMzMjdva8bDfB4/AEil9M/LIOMb/
pTj41BWEiVzR+ttnj8UQXf0zFCixA/Y/SE6ePDXHvEig/2Ap9N8OtGfzhL0gl8kbA6Dthuulfj37
cRpgiLXfmnOY/OdqziMtuWupHcYBhAnz/bWWN8hLRo1sSiGNWCJV/ATUzy9bt1zGskwaIx2iKEnu
ehsguuGimfhhoUao0YFgoNHeVjTzTacPpyj1NHPgfgziIApdFu6q10JvhRNHR781FlJuv1/2NwOw
lnSLigte93hm7SMODyKEfSnQ4VUuDayd4YyOp/M+qWv/iei/CbiIFpzaDSqQZfsvHwl2RWGxXz1U
vBP4/VSkA9YyXaOZQKRVmz1An6siNXXZWchKYKhjvW5ovqSBMG+jtsKKrrOfomJIgoYcUDSYE9ns
YNN3l1XKIf1wFK1Ph5Kg3ODTEuKy/Kan88yskeZRENplMhYi9Kj3w+DdRXfyGDJjfisOj3j4+cKu
STgGi4H9K7bLkpDvJHZydyUY4ubB2XpymREzilKHPqwtZYc9ECqcP0dsOUM2k/1skc7i4g94Dsaj
u4vyiPUEX95gypdMSGTGtRsvtC/jdm+bMCAmgNxpx1UCqx5IucDFhWLuC1ITKCtt2L5ifqRf1uAf
lQHTEYrEu1kxtYMKAvPIGX6XMl14NJZBEchr+sB+JZOC2FkUJNbI4U4xnzZMz0KPShaUPgWzGiOC
x0vUrlmbwH5W+g7Q/bdYMsjG2jVL6/kxk9oxWFqNOLJVH8PqqEnc0+GTFWD+QAxGkWaY7aHrRw8t
tqcHnuZ0HlHqMMs5gnsmuQXMecMHHk3pdY6jpx9kD5l8wKRxFDvo5c2o9r8s8MYCWX1RzRIKZR2j
Sw/yD8mss4hi/XOD3brmVzSYx8TewNzNzBaXej47cBbxqPro8qQaIG51u3E2Sp2DIer3FnQgf3qC
dlJvLrRGGeGLAbnQSPWjjA9ft+vRRa6m+NXdPdLGT7oBFKvSiTnSPJ1ybl3zT4mW43YcaX2CX8xe
z2YdI08zX6TTbrxYD5kYjIuUjdnosRkEQzVb7ot6sAHCGYWEYDJfZHP+kkSunfxI4vMBWkDjQDMs
JcJK8JQa9Fyvxpbq7kGd3LwITVwrSJHYDnB8a5v1cWlud76e6GB4A7FZzSTuoAt9qRI6pxDfhfri
BAQGE7t01msaoIjSNbCdmTlEbXDsu4wxodnCRcsfkZ0jGwn2Lt5NKH2WNSLK2cvu56Vfy1Hn76i6
YJbL4okMJ3qVd1FTSiBtxJUn7isUWNlCqYvvImzhjN5foZioH2/fT/P9IzeGgfGG84F9MkjdJYnq
IZomJC6BDyQXRaRw4oFDj7/LY+DL+6JR3smeRz1zHza2knZwbMIVqj0WFde81+lf3YQHVzvXu0/x
faLTNlUccEThETz9Bz5dc+BpO6iPENjqwtL7Z77uYrFIdDFAJxDeGz0YMvyxsNZOUHKoxN78VHVf
TwxCff7czqFi2L9lunMQfr4k8ALtEQFCwmMXEOT5wwY0YII6MIbyhkPYRVyP1+dz4Q5O65NM/l9B
uABc49lK3gdTsoxosnOCVf0dpSDuCfIoWaIx4pYMXMXCWJRt9Eq0Sj5rWXwubO2aBCU9SfL6z+FL
9VR1NLKK1TEoORt3iyw1vAAajQ/56RGEU1FPqVswFS9Ou+APh3xf4nAluqYNxZbCZub6Fzv2XLLV
hImCuhNf3OS0w4OVEDhx7YCrTFZLSQk8G/5E0SNK069BQQsbo6DlpM6yy+lIeBq8EOc13urQduwL
YnaUKCmpo1s9HNm9+ZEu5/y2HDdeBcvdV9BNF2SEwa0S5T/PaGm16SK0vRGiSMz6HX24NeX/pNzp
iKwee96BLBm+XYWni9CErdlaY+RUauE8v8/ZhzmIdbGYLUpUShYD9Oew6VTVXw8GKpMfMMNJiNuK
md4mjPkGQBwKhdMAV+PYGwXl3h+rFhhhErLLBD4+8GSrnwdicsBqxwvMe+s+lVvLGQW1LVXLRvQj
CyTdFm6KmoKVRd/42A4PjDH+dHChlz7cZhV3YvZJiLSdcCKlzele1EhCC//xr6HbVZO/Y5C5NiKG
g9LKA2sPZ7WL4ZD/2NSPkKBrIivNOAJkFXZfrpM3a8Ar5sQEv5/zZdA3teLDmqueutXTcKETDj+k
pFQFqRIpNolnlMrFtbaqIr0YD3AtGm3hfiA2geZdH+xzctPPUU4N2wOXB/wk7WdgD+cemC1hy/eu
0AUj+JcNqgUZHTmZ2mu11FsQOy9cVOPL2MwDQ3n1o3rEBsrLdMDW2f3IfDEiQEiyjYQQpYSFhLiR
6R/FNIF96bQJ3aNa0eg935zQ/GGwTi8KCHuN//Ih08hYygtmz/vpKBtz4eXd32FbXvLRXSAhQQGe
CkPyNB11ykOpui2PEKDLQQUUmUJsqUZwWY+2V0Mkxyo+TSyWYWgLO2dYSIGUIyP5/KNyrek3IXZj
eaU+bBKg7uE1ueVdc7RIaLlcUqJugvvCiyqqgBxHBve0S6AHA6MeDRmySAGqlz5B/E0LF37Cwapp
mbq2sbjEX2waQeqkrLeGtSDG/I1vKkcW29zDmRdPX6NXzOQ0w3ATsQV0Yg+X3S7I/eLJAYLhm/uV
kWgC5h9KM8Q8d1X+Gd5A9WWZl10FaoG6WZqjJvCYa47k7Cf5cfTc1+tijTST7LlnJEVBJTX5MR96
kbx8YVBZgnHfbvjEkZs8m0Y3NfiwJMHsq9S+lXFsXhGidd2c478VWlo4ukFenTzebwLZxqJfIkuR
04KvJklHFGItUEjSxi00PBYHa2XX8UIiIf0UjJ6qqDUYdkJB8sJy2vqGkVuhw7c9j5dtvsru0h41
zymJ+L5/69u3aosjh0dSmdJ6wIbDJHMRLjMTEc7PxhGbTpj5JBolcnyjj3+EeM9KItQTZb7YYUqh
XIZW7VEDh/GYIR53PkhHmj6ECS6pEVHvZg6CgQMKFGFKekdb/ZJg9kL+SztqTW27ir6JfVzy/lZX
QahTXXy4ci59M8fkTxNY/NxO/4t/Dc8axPQB4fuTum8ZWd41cFUULew4vyksUw0zGLrtYma9eEq1
8pZeNrOG0diHR7C+80dlDKHx7Rx9Y0NP3pmJfnLehWIURggbk0a0GtK5g30NXHtUAGVhVasGygfM
pf3zmiAeR8OHaGRbyRYCSvyl+/9+Almp+IwpobnN+SPTZcMmJPixuiy0aastDNeJmvzm5OshUM+I
RVrPeaNy2Fkuhi63BXmuGtJ//raAwfDpN+8XqJQQhIabDf6W36Hnu8uVJszxEi0c4a9RLWs7R1r7
pFtFGvLtJdM91g5Sf0XP3PT6ydJhnoWYNRYcjg9/r/MXrhkaCcUac4yPctFQ5T8t9Wa7X+mIl2xo
2MQtXmo2wJEVpXQyYcst6yhhuFDq9QyB891g2PBX3YNL9rRBKwOhbxa1Kyz61WsnSp9whfqV0nfO
3/G9jTb1/QuOHjdaGLAaSZVXiCw5/+ahFYsU615Xin7f6ouosxBihIEPOn3dOm2sfgqjdN/aRXF+
q0GppQDpVHXzzA24HObbIVQM54BGNTI0ltgXJvJSRI+w/i1w8kj+7StyU6IV6ZbaQ7F7uSrTYTry
xpHcsrydD9/vywJtd3gx0ank21nkAuB2/og54lXLsQdyasAI5++A4jOWPNPBoWcMzk3aBnATAo+/
gHavdnxIvOfqeE3Q9zvmOnD7FK8r1jA5PNAI06D9PNM+NSlZ73RnTylXzI75+wQQrbxtiC08OutE
b7gOU7fB2upjnE7sXPG5JQpxqd8s/eXurYq9yt+rWQCqJ01vIndXHS9DWt98kN//U5hYLQhS/5fv
bI6u8YUbB3Glw8x0rPhhfgK3UHZ6OxL3V+22sX5Myd22xEPn0y3BEDy4BrWMEK/Fn2dBZqedgSYM
6c1A8EaRi2DuvWPNSpG32MkHCsLl2zfKR0nJiZhEVMzRnAh0Nd3Zb5Ix5hiq7OlImqmD30zLObIi
3G+DVGhSNgupY4XLZN/xkLqHhY2nc3r/n833+Vx3oX9h/SaSPJnA+9vRs9WI0Yl+FY5UEqLomTew
sCLLAwCkBxhXR2Otg/hBycMvDWO5k9HZs6NMhtSizGbKG06ysJSLr0pqjcHcCMpKwxSJ9yJC8e2Y
8WKog1ld+zTspUp40Nh35PU3SvT1Rv3oahIK1u8JPgTm1PNiD52AGOb4XRswZMLk2YhDkHxLs1/t
PG89uMN9uHll2drWqvtQqJb53XAzt0v1XEXR2X/fdasajaaFcozvQluQuaSuooa9adrkNus2hhWx
JDZR+bh2Fk15bljzYriYtZJILhNDNMt/IlK6RJN6eH/gjGJg+FLEUY07DPxmLQ7PhRY5UtPeWzti
PhntF9KEx899ofijVvimycjvjEEPcWTdVI3NovNay+Sf/+QvfLco+eVPCFSGFFRxaVCtSYKODgrH
KmRPYjdfUqY9jKESANnCBGrKz4Blx46cnAwkZeMG2J5eXbZhjhHRJ3LblxdB7DoEBWPyPJAPeLau
vCwgLW3odR2pCRJ36yZg1nOMJqkXRU0zxs3t8fX4nd03kBS6NzxhC5bDleYiEn6ivEcREm+LC/z+
ca0Gc2/2SmX/QAq2cPCmKtA0CPvh5g41DLKp+dNI+C4aocEieztBjeNSgvsKvSAxwibhfppgQs0G
T7AVDi7Nu1DUu4c2dr2Oce/fWqlJRrjCjpIlMYO1Oxk/G1CLcD32cBibRhNa1SNhKpXZ12F4nkgU
StpxFxKxPMsVCvVaa1vn2bt1Bz6V3Tag2bqgX2b+gNBvjR+97wkjXPTpM5Uh01kDqZVy8qM4S29Y
Z8a8newyoJhjg0rC7XrrB/jPAqSPmESWa6rw4FCV3VWEaPNXvtTPX1rttI+hPPZLuzJXChev8FcY
8FB5CAlnhGQxJszjpPkVWlftriARujrcSW9hS1ilKvt/21wyVS7xOulGb6mo+/btdgixMKAKJ81s
HK5rhtgMzsGYkmAn/JdLlOjmv9aYZO0buKzMzh4yGY74P13gx4TvAT9vPbyayb4CXorW2qHDFAu+
mUdfYc0Obu/OCjnsM9cNGBiTFqvPlUUfrpxiCRm5fwxxLYNhPYVadxLufWRicYDhcC2/yRP1iBBH
LePyqeqmSpBwo5Q+0v9gnIObPrZ+S+gef/Whn00L3coBgjG140CpXFr48/4l9nnXbomiPzGdXzq2
XrvUJ3DgH5bBWY0Q9P3SbRA872kwyWPIo6SF3d0px77nMl5t60fRkSyr5eF2r79WZdDFA+SCdaVk
xURbF0ZsJ1gPeVOC3bghir6iJva7PJ1IoAF3a6bJR0elXxLuHsaAEvjMs6vskenCtrYp4qEr/1gZ
c6oMBw+Cipoh5ECuSpT/kQwF3I0DN2oLS17rdqwXFtlc04hMdI5Fc/Lvp2YN5F+t5nUdaF/F2JKi
gIt3z+E2hLnN4IVzOhyit5FQDSWolLtRFQdfh0cfs3McjPeLnvtUA+CYQiM1BB1Q3DEoWbGfC8m3
o0wqyfyCPuHClS2FjycbIrLPZit279TOKnAg0uuwDmlMWngbZ2j+UvYSp7u8zyTBgyucgTtndIdJ
SUFeDsCa5z9BDZFMlg+MyHUMry16mD+UXc3HSxDSvRDoAA7sllTYv4bEmMOlRErr09KRelKGrgwS
v1L9Lg9+XjchFN3/4Up2/44sAWtwze5QAjI1ubPjYsM+GwtCfeWx7BWTfDsxqxJpqQxdMXKTQ7n2
DrbUN89urYdAKS48AF8TBlgQC11XIggER3OPGhb/3Rg3oORyieYYaifLRKZl99sss1RreM5/F4A+
pL7Quvd7nQr/rJ4IdoMTMhd+C+iqjLo9R06TYbr6uoDm/akXNAK4v+iJfDD5q3GWbwp+4gkmAwce
AFyjVMd8/qm/Gq3jkGjY2KdWC2SSPAPXXuzkkpWbQ1lb4lvsiORWI3tNCJ7pNl1QYwgg96G028q1
pNGJlveuaGQlMc60Xz3ICsTWxlO+Sbet8udFPRIPoQ8gIFBMT4TuyEx1/CX15bkssiHqgHTg+95/
jJP4YTn/jHqCW5RlYC+IhYfISMzSSnh1HAtq4Ab5zWSJ1cHkAOob9EIJkP6J4Pd//sciN2RwyZU2
j61ichRTHPoQnekR89nyLRkb2twOqg/2kWF+yUiruVQLmR+uAz4QmhGzjrrKKBzD7zCdO2KFCjzz
mOF3i+H31Y9SnWGW1x8W1ehaKAssD3NcfJQCbAwbdq75gohqtyhp/MdPnOGWMoZsv2sSJFKswt5H
wgFIZSZbzdt0euIDkbUGysX6esF/KqfJeyKfVDb2s2I1K12Mh0D8A1Jeg6wxhtvdu5ahvTdPIm9L
cwHSWrBLF4aEEgnd/mJ/hxm0oKuLKK6rMGNrI2o25wTSlbpHechJR5Dlr3waJk7Ri7Tp2/K49of1
S54mDM5yI3bnqr6tB/dCkDVSeDeBEy2LJNb0S0K7UpkpXwKyMYKxKdZ8A6pApkPYhgu1XYSPKnbX
J5JSMG0cRkfQkRMDT7u8HJNJKTmCNp1lWy/BkUALaU5UyPaT8zyipUSn0vUNFWjXi0A44U9MFQg9
YkFJjc0Au76oI51sUfqPFNhy8UBMdGjDcHUZAPAec60jb2bzHESPRa5wy72ORlM61s2kok5G3TOd
B09jRqekI9Tmzs5O00VNzx375y7fwJOk8vuIhPED70mvTX9UqldAM+XNR18jtgfkNzXNbqUKhN/u
rfJEI745rqMH80rmLi8DnQuI5SJY/TtggOZhYzbRJZtSwOM8n/CVmimX/P81+Ydq6RRRuzgjUh6e
G9JYMamJgxzR6pb4JWkNIa+9ovRgUPPtGFZzDHSE/IWq+r4m4TWPRP6iMKWE/IoeQBp1RawJY8W3
mGJ9duYIBOd1ycZAA2mq/r7ak7EEYV5aWFW8xydWsC8uPTAKy/h+JTxnkPPcmo0EFayqdhh7tCEY
dXe7T4/obxl3pCGib93pdD6zJ9LkC+C02+a/bYootxgJHHTIwVrUWTS9Fcdqdvr8VQGaQQ0qAAbv
tFvqjDO/KkA8tT5G6H4TqfAMvdrFGZKu52yoj2IkjZT93RECU3zmfrRZyLG4KVOPjLTOQhkpXdcs
p3IZiLgzDxRloWqek9R2RBl30N6SSVqg0K80SUhYMNjvp2v7NpS9aIzNJoTzgTLKVgbr64BcVwOi
fVU0MXauqQe5iG3DT+v7RCsD2PzUJYSTXz3c0Bt1KOcSzMw6J6O7N4NZNtLyuql/wNmBHCv4s7Nu
UWe//279M07nodU5sjs5MqhxtW/lng/iqxqOLOG66l/69lyaoK62WetJ8xiPdRwNqlCyWQeWavoT
FUPq1LPqYsUUnAnI+XO3TFterQRvlhs0ttMwTcBAmIjUuWOYqep5L5MKJpixjHJ0rMVziz2N4XFy
SmPrIgvR/+MrEHZmsNKA71rMrnpby2ITbypyE487eCRtl6jwKXKVKJTLg1w2yQ+3z3fysLB7SOE8
mwbh5nnd5xYwCI4UhAxvsrUcPgsFrkIewz4hf/6PFUcl2g97HWvbm6uQpFTjz61XesK4iVy+qBAC
F7bh6nfW/VNMgk6QbkJjepfBljyBi8sll8YBcWRWM60PeT6kMhvBibazhkIsr9A57NxfnJ3w9huW
UmhFFKEor62keTiH3pUfPchawiTzCzh5BblgZRA7NgoOVTDbDXqkf7OZof8EoEFDMTvaOO/DCOSo
0JXPj/QAdoqrM0nasqIS+Tz4/GhqbH+SQIQ/vU1JIbrWNykj1kerljsUG0++NvZU7mmdG4I4Ka2c
2Z5slRQq3T76n2UhowrVpzmiFKaGgOcLCE3uQkm0bC2e9oSDQuReddc4Xy5ZKqIYH41bEeeZWkht
VbQDE5UkY6VbhgY6Ph0/EecxswrzFoYD8UX2Vsi7VpwI2xMPKtIbPbQQ34tXfA9N/vTc+r+S08c1
tQKGO2NAcHFmd/o3k7LOH1+g8Qd8/SxTQV73t4124X0HCHHwPiHnmDAr/Mpe26k3cA/iTfR8BRwP
ATMGq3rnmbl54Aay/rS3M13ayJNXC0CfDIK5clhks6GpA+O52ox/1jkF8GNZ2EuXCDL3JeZhLX6T
sDu8sslbkE5wjf8wDGooKDAH3vk17aMcbexdDHSFJ3s6p6hxzUoWwM5Dh+1TfnNtix7II3012Umx
8G/t4yMV6E0+xrIAUcsIoMV6k1PMhY5TOyjDzCQ6BjymNEqsrB8dC+cxI7J//33ZH3dbtE8R9Xv/
+Xwvhqp6thwIstoF8xaARbFYTxk6a90F8isIr3yXFgmHLZIa0LsS0I5zohkSpOiCj5zC//zMV6f5
PSDSBL7g+6Rn7e+5WhW3ciY7U/pQm082bYUMOXzm0qeByBvHg8wqmAqB7UrTCLFUGZzJzM0Ftymy
jM+mjFek6cWwymiUv0j9jQn+xDuxZTQKYRDPZm/11/vFerwA+/UzYAsqnpvR+Te92ptA4y4HOoxJ
+mqE3dovBOjFOE5frHI6RSo73hMjvsVNUwPOEbqA2CXcUhR0ta6t7ynkF+M+QbYzwxg1odVcsJQ8
FH8PCUSy6JgsBWL7HcS6/tv5CYZBNpPS4rMPvF2gP7r4awKJld347pkGy/OR6dWsf76F3Uu2DUVd
OyG3Wk0LlYExPdw11Td8Pn+sjCXC5aYSkF2LheE1QzsM0/fQ7crhmZfDTIB9tm1cgId7NdGX2DfQ
CtS6ONLw85LnNsLgT8di470vSQX6Q+sBI7E5Wc3Ik45ptrj0VqvGoXEUn/mF8llKS4E25qw2mHNd
b4eSCX3DaCRKOJdwgLS2/xezhkmBflS5cXS5JHYjMkP6dNiAgRFfHzg9mmEog8pum9GSSkpG6TKN
89lEwbkH8JZ5+PF+QbAYC3Qw9LxphgBKirsYEJpKUxK/ZUaa7SL7iKP3JSIdwmTA4KyMoZy8PkRR
IGjH7bgSFRO0SfkagfmBJAhRcFT12UeEyl+uKH70z10MEl0GfFCmbu8nc1YDokr0y9RpWvLRg3v5
Tfn8ZJq4qd7p8bKRkXrEc4fM99y6/TfoPpJmluv4RijABB/II/ASdzka/0mi5t50OR0Hc78Q4d1i
VWhAUl8uIu4qkGjlOfAkgghkq+QcNxP0/xFIgIYXRCwwMv5LEm/yfZxVhsY+nxL5aR0lWPb7Nh8P
rN+EleJyPbIjkxXYSKOe+5ch2Eb5EC3KpoIXviraCyIcLhEM8tgzYe/8971NnyVf9xvIgkeKvSLw
6ha2+4sriK084zEhz6V6ridNl6QTyrwBwJXrJq2Hz/gP3dkvgyhvzZhgMEOCpigwGGftYD+o3tz+
DUvneClWhL1MGL+A1iMN9t6qVZ/J3DFkDqYcMUqbIeRbTlCUYjsyQcR6XhkPPD7eQFnC4PUNxuNV
5bAJoJSSsV/c7U7c3oKK9Laop31x8cULtPTTM9vgqv76m8MOvjLwciIK6tk6PhsdQtqCdlEwA+DP
VaMdJQUJRGveUhV8a+LoL9Ma4atpZcS98yQUNMOAOwlljInW1639PWwWNAOonOQLAhfPGZpgDy8H
cg3glCaQDOgj+fGIQNHFxbWYVYerVT8fpazGiV+zcnINOa7QBp0c1I287KUoz14RaAG02J8l6bB1
O5rnjZeHnAz5utiUAl7LT1DUOrspFipv5p9uvYO99l7hW9LH/Of3Isame4/NgLpVILMKyb/xI64G
8j7YHMu8AsQK261THgXAmNn0m7mzrMYWummNHjciMsfAKBOPsNrdJpqYtOyLGAWOMNOysBedqA/k
TteBfPEt4aGuOiOnpVwxGS2Sox2OGPiiZ12Ad2Avux1y9/V7UtUI80UsRQxziFhFd9brc0dPlEcT
n6D82IwdY0L+M8ylq11F1/6QeTaRwXQncQrLmlAhyecBtIFPaZ7Ca7SQUIqPz2H54xP1ia7QdBNA
/kd+f5rbSx2/2Nk2dLDJymOEe8Jtk9Dwf1Z4BlADSpu2Dq17Nk0w/rGG6+Fpyo/7rFnjyecC0Ll5
CfhV9lCQqC3xBI/jGq3A10xYxT/FYa81IUsPiifpmPhKiK/xhDB9w1dJG0DMLMWGuM39yMI5pcIy
T8K5dG2ZYFBvH28Oc5CnldNFwdaAXhejWoVMzSbRztEoBkcWDhM5fZa2vpZkVS3z3yefFUcxPwfV
ngZE4fX/XPcIWPAv3MP8IQUbuzKGvDPXpL74qMObOm+iijAYIbDYV1e1niQKlw4FdJulQa/82pws
1SG3lse3SRFThaO42oOmFTd2DRz+kIdtNi3dNAzQRH6YzOdqsLg/9Rxp3bHTznnpOPwqTtDAibJ7
gLAwKXoT4vqKv5gK+PCN0+wrjF/KgvIHt+Jtnw8AyJn4i/qPDrQZRiUCl0pnVJDe7N7EkYAzOb/f
lK0Cg208M4uX/Itkbn9hFNNUOiwPIpe+Ma7ooarofpHubQkzIlj35qGW0ypPuu5NHF0lEvkf/1Af
UHG6Ql/vT+3K83gtPrNsygTP4rT03Y8dMoIorMZZVlHSZD/VNVCnqS/NkRNZ27Od7okDrTzjz36D
yaHi1+dQW1pOTfBt+AL1vTmGmXvtRHQ+PMLQeE39iMPNX9hr6fjz7l7tIRfaDkslTyjQHD19r+B/
ZQiEYZ6H5JjxS+AG9a5CdWkCFOhsCunoUddwBv5FoyJ28dG5OtztOugG0pXAGuunZFZG7TGyJkTc
L2LSU5huiH+xZsdOFDbuOGMQ8wlk4YcVu3Xy6cYMKjTm5b+wTWbQed3ZQmDa/EwaEl8UdnZCHI/E
YdepFgZF3/n6ST6mSaGs78WYyy3T+Pj8kpsKkx1qoih9n5rgDyQW7ibArEgTW+LjeE+HbDfDek3S
TnxstFyyQkrHD8yzaW6bTOKUf/iq82TS6ZXAIeQqAKn9OBuE5ap8FQc9GgKI2T415VRBUddGRW3n
DLox+kuuC2pTKUC/33ZeRTWxZOe5QFr+NEapsfy1GZyuGDz2qU8BmSGmh5+x74SNUTy1sRzP3kHn
odJ7pOddcHnzdfQbS55+jBaOmAhbY1RniInWfM1Rv01djurcJL0BWD81KU0OF47zyGSdSihJnEtt
XM6sHUZ8bG94sRpfETw6MZ4GJ+TNjw1hHzjf7Zm6YO46x7yz7lPn5zLAC66kB94xkJJh+kIpT2nB
P6sS5kU/9awCJsl4pMmdZNyhCtKofXuRbdv0RbTZeQbJ0E+j5eSklHYfQQPP9FcL0aFHCP4r8K3e
Gsf699DzVPAPNESPiMrUDXCOgRNGh2kh2T5a7lKrOtYaiSNIOqJZ8aJz+VWtBfW9WShRITUcVCce
m8zrzf5cAr9UiLMG2Ru9gm2RHYAZmelh3MVOy5azjPTvhH1u4HhaZtpSKODqftvKg3ksoF/jPWYD
TKx0ZohpiDazGAaoP57MDrTWK703syipYcl1iAJUfsEPxS8wHHZHw0yl6h7fyXQ11JKVXHBG8Jju
X+5I5hzYxitBgcPb8+T73AaIW5alWhrbB3tONgw2LNssdXBajnB18inFZtia8UsmH+drxOxfQZM4
6Zdsm5gn6LsJdZMiLVZ6SoriKEZ6zkq0EMMNpwE9VAVU4Y8QTslgtXsdxeOJuWFoKhFcHpDyrmZR
/XGG3/FOHHxyelcTfdVbL/lV+BKUg5ilBbXa2EmOtBfmhBe5v45OfT8dePOV0bnVRMHyYU1a0FAF
LQl2yNDU4sYfiziEgouxZ5HzaydUk+OC6OrIW8CH1b5fyezr1lpFDd5UFm6ZhbdgAH91KsJWVdGQ
G6tgSWDmOtqReXZVYyDoWDqdY5ZKYmrsY/SrZzmQRm/ndsNpt/ykUW3WvivzbdDATq2bKqZPSSBG
fBV9XffqFMqgSvA5KXn55HYkRhr6y2R9eytNl1oco2JWLhVaY1eZyJBoSsL/ySnmgkZvsifW8anx
r1PCxZDZ6j6MtEsPgvZzY10mXLzv/DlHJjvUoxsGdoKsc8sYdKB8jH7O3vNQEDM1EOMnKN2SQrA5
8I0yDUXBFi/DnsSA6RyoF+U48w3ErR4AK4evmt9+Jc7llZTS1lYltTVBQ31YnF24cIV82mgz0o/f
f3iX0gbAqmZ9LDx4oE09eynZpDvWwrOPnxl0PpUBulqAw9HDtgJ3yI4YWuu3eisWUXIo3xdKKBcJ
KlIl3I67fiLaiix6VM4C+x6JwxS2n2wBosjchAei3/PJ7qHkvGbful+x1ysLep3z77kRJXVcvxf+
MDWgscqdJ1TtHzEqAxRbQgFRIaI1P091O+H43Ddd8EqoO+NYr371+oMRzJYydeqYAxS6N6tS2ihu
KG8kofBJloLmx97eoR0khB3tWOMbMq8fHYp8Sz4VEy/KBz/zGP70yNUMMX44+RBv+Lm5d3ShPSGc
n8THUc2iNCQi/A8swH5Qa6b3Bh207kDt2VrHA1s1emViACNBl8zVbAJKno4dAj4mmiN8rw4iSulD
yPLBdgywsas1oST5bBntJ2i0VbENj3krHM5Jc8Wv1f7IsNhkGnX4Jv2Jp3nmzetuuOU8uG8upX2c
fh98UjZvhMYzSDJ9vx4B2k7+DtC0kWge/3ddMAMJrM1iNvjeKEerdYI4pPahC0NSfGt8C0bPPxeJ
GyGBC5Rs2yXCWpdzpLb9uvCLhlHx6BlxWgQjevk6Ij+jFjvWA+7mnqPRcNJtfy2gTGqmdx8Bc4Yg
HeiDUGfBZI9t3DPw/Ti+0THIoLmgLfWnSdiqs7y9+1Gy5qtNRFGu26WSy2yxFhmJjgEcHUcHjd1s
dHsCfvEwo3nCTkEuenPMBggWB5sNxA3JO7hjGoEJug+hixNl+WVm1YLDP3wze59Lf11eOwDlvZra
y4i6X2ZgnQEbkwoQRC6aRuSAa+MBIMA7QXmczGlP0jYbXW9Rb3wWIfOGiIvOneKjb1UXm2S+LlQM
apAigi2NlFWJdsG8Rp/ZPXSRXUQLqo2bgOe7vS0pC8JYcVVIrmbZq8zQVs6w7BAGqp2tOKLQ7LVl
5BerlbsLpofPPfE32X24Zmb/EKkB7vq2eCfrZP8DbFAeKxVFf/n6OHrN/tfuvk/WNlhbDbexANjn
n3zcrF8L+G6WNX3+YJy++V/NwreOuwcGTTdkkjQbHOT+iapTkOjKg+fWbLmcS59/sEKWgJv9S5TG
AXbfWX0MPod5fNE9yGwNtQluabEdXMOfeoRwQnoowWwi+cRdiN3HrHcEQjVEIDShvjdk593sDMUn
FDL6oZJqpFmOYBZqH0iyogSBi3Imhh8ICEyDKlHS8r0Pf6wul/11my7CSHL5P7oo/3wHTy2X242L
aKN1ZHwKy9XlqD3RVrEaTf7rnSsU+sm+ad961BZSef1TyEoojSkO+MtXQPc8lX22HEn32WjzlDlH
Hm7PJ6vufbJ/ZKra3HsWmChvwPoY8jTJbAZfSte9TD5jH4+76k4l17Tl28kvU0gibgSrI/xuIRch
avTDz67c8EOY6wkUiL6He4n4yqK3gvtmQdQ4U+X1gJfmnJTjnLhI7Hutqejiydg+fRa2U9FVsarU
g54CGi+1cUQzr7PFGyUSlPDz4Ey8hBftWG2/tpdvJKXr1/Cn2t+8wNEgGAuNd2LKoz0Ac00B5MjT
phDhZYOVvVZtyShKUQtiKU8l/CqQ4M2LOkWqkHPEH4bhr5VXj8R5qcHk1tTP5A/V97nGkqtE3QDh
aS2XV0d8tWGOK04aVrQd53ll94EmFdxoit6p1gkFHqaqBLV836xsMrhnB8b8Wh2DkJbZYGOeTfXL
jrtGelWrF+34Yg9Ub2MmWRWK49OtUGye++dnBkkVoU4K5EFZczVyBN6EBCT4j7tCwd+HvJCN/kYz
tQyI9QE3oXhTwqB6nZOhWZDEfRfqs0uXlp1Bob0b7bnVcTiV0q5uhLy9bkbWeltatZi+JBbfy+MI
rriRRjM+S/s2Thd3QB32TawcFxZJZaGM1vuJelBinK6SkHa1/VYBHbbjZuhpKBUgpguVjWXhu1e2
QQlBbz5wdN+BhkRV8ZUEjkDmqYB+OIXzPT2Mr+tMcDaadDFCTbnogg6jXi7zDmQWAayI6tQgq47H
NppbNN9C9lpdsim+GVnF/si4JvwFZ6qqP5W9T5Ko1+M7UQdUCMflXe49msponJ+aWZwV83734r0+
WPaX1bRLZVbcwKIch2sMqDZyZyU9MR5SR/iRMg5w7J2pfpRp0jseaaI6sBfw6RHgXBNBb6w9QmbW
9jhpOxAk2UhT42HFnmNGj/X9J/n4AMaxPwZuYRzLO8NJ1P+/37mnvjtUTJw0j/uJJ0+Kl1zlMHrO
IEtnj1tPyKiaPDrjXIanARZFt9lQ4XTbdthC3yBoUjT8WAuYQBcbJ8LV1oK6S1EhepwkjAbSX/iQ
ZEyDhWRkmG5XozUGWUJ+b3TMzkMuL7FjAMYJ0sHnIAajtoPa+uBs41bPitrxi7mGg0flJklcMtju
XqacATarpuSYop6riZibO98a0qrkjO1gxEamPmQOl0WV4v0laTlSD4uUfJxyIbhConTlzzR1YWQD
O4byzr0xQ285BeJrkUpfUDV61FCFPmybirfBpaKatuc2Umwj0Bx3hlmVWr3eeByS7ONiXtHwmWyM
3UMGFRgu2MXxZEAQ+1urxhQSoPMe+1FJfkkQE/czpw+5k4rEHPUhOIvBrihORWzqHI9zpJ7l0Liy
fn0yNJXl47EgHcv0FBtWU2PZ9xDHTNyAZwV/4+akNf5VZH+y1mItqtHvUNyj0GcJtcSyCSwBf2b6
WLN0Pm3XuGbn3MW0aPtjvfxonF5qZifpiY0iIYL8VsFcHGEVao1e8SFHB2KemlM3NBDCLRUlxnB6
LynxmjbSr7hnuurtYndKv4FJWFU2LwWrbQQlc7wBOf1/ywTT0dfvK8pBGzRiy21yQ5pRnnMkl8df
RX2lb31Buxg5NT6auASH4uOI8z0ofEOWC/M5EIHx6fdfgCBtbhL63TXw71ZcQl74WXxBp5i4emnu
3nPz3t7Mqxz2Ywjw+df40LD8cGxCj7LrhCTxSTl8Pcle3282DnQwugvlQf3pi46wPCm63JdyxWv0
n3G4jZ/5NBDWMI+ZE+dkcEDGfK48hNgheUuPeiAA8F6PVHxOCeDAZaJ7Taty9y7Suma4Zn02j5vZ
tj7plDg6KbsP/WA4HgArW7OVnps0XYkdxtyttHX1gYgycrU2lo5brMpwDNn2LcMZkov19lDGxUrR
dmJutVSdDP5mNkdZfTRhMHGPwgppGGWdMz0VCxg65tApMB5rskYb55lhVb/JJCvRoq0UJwEZTa7M
aLNDS2Me4KBszJeLpdTZqmUpZT1O7y7FkBXVYnC/fQ+DWOSAhOKQx8Gu/bdfrtO48yYlbVh3KLRG
bZrwSG3oyREn+fAizwJJAc3BfkKodvU+UyPWH7mN7Itgb34jAZHStiwtZb+nWshpUGdrCbPiS7+T
Uh6LPuxUJNhHvId7A/4E4GfUwG0dIaypqdwfrSaLTp45ql7vqR/Az/PpVYS4dwaUEBX7ZM6++4Mg
4khichjFLKkYMnzmAZjFNKo2cWwidqML8+R5HrHGnllJDwf3X9D/yyDuEmyiPwKN4/EQxkHJrowE
XJiVlXczdP8p9ezuIzeDi0Umx5VfZ9rHQU8ytFGdVjDCqcPrANM2CvckRtFCzJRcIjVTr/iYaWTi
eMaaZVzAT7oBYUcM96z0JMfxpDIJkSNPMWVzRX71Ez25ni+HoyEGX84Q24l9eQ/I0y+N2e5q1QPi
/E8QqIUtGgiEFO4XYqapO7IyJckh3DHqMMO6iQBQyyaNJuH1CeMfxNw8iC1OwVb6hgoHd50L+YNm
X5e77b9L0nQ8ESRG0pfFczW7n2uu8t+z+olcQOqqr2LKtBQPbC47v6NyxerI8dIKrMZh0N2p/h80
FXV9OQPdeWTh3SAll4/TyRSGnilhPR1fwe16f4WM69VUf6K+l39JtKstoagKkcXDKdyX90yHhkPR
B/Vrz0jDg2t0ihBHsvLkjESUPp6sTDu/xlm0BKn8EkmpnngekkerEu3AYoUwQVcgs28gqJVKdxF5
FQKTBLp1OOdOZ6rlPX6I5YtE1+X9uODlBMyr72LgVnRwt4ROztG272E+MMApssmd/H3+feAHVCHL
Piv52KFjCcdQcDVCWFZlXlj+d8y/BpwZuQZdSqUTl7UDDq9FiUIa87JHZY3DBApbcm/riBXD5doQ
XaeSvhhvBsuxgSw+dC5uGuBKx4WCcq4mzh4sk9VfNE/8lXBIP1rOq3NcHykRs3SxNu5XlmnHA5pn
trZ+TOhfwL1Ziyq/O2i4kKTJr65rJxe1RWBEwwFCR9Jmx0L6j2lHmJ5GlUU0nxMDwGcv9HSARHEi
aBAl26czuPZW6J/4+tlnNT/l09WTW/qx2KCgUWAvVYVpaEZi8ls/EH3hJ1450CJDSD7goAaKor/m
t23KgPQGRnVjE0NFRjQMNXFdm7Ew3L1a3FAiU0gPl510LYeVjr/NevHxRERKTJ9VaGsrfUxjG7++
UNI8O0Doj0AhIFUBV/zhWmUj/JSR68E1Nftep/kOENE0ULhb2kd5RBGwuIYwhWok8aQT97E+8ykR
y9/XJCrguxEAkGeh0nDVpfoZALMHlOrjNKHlnS3gexC9xqIURnXkgIutyxP0jYlm37/4BMaqcO6e
wHgUro0nXSkdJH6bPRU/tVOxLvFx83YjfjoSJYP7VIlT9rwae97yPCdxhnIc+9AZhY8TLw/3SH2v
LhDOv9BEoF/LgtXBRsETfttf5mUx1tx6Mc9G2DmTmzM3FgG3dAK++lfPFHVKiUSCMsUQi+RnZh8U
3Y/JYDOvGl4l1jyttVNMX4OfKgYjg6hEUTYuXeiDMOuKMAEWImNx5xEdmeQM0RwE6/LpLzri8xzu
UL6rjP1FSYGf0dOt0LMAplWPT29VjR/krBTT2WFnToueSvdTBTWFm1tEtZzU+gUSWFnGl0d1wtkM
MiS6wdSXcJ+kmBhhEVMcqo+KQ2XxPM0XgzgKYXWsjIxRcoLpiOFznibmBgd3qbeCcIUvPlQIQZTw
aza5c8djQUdKZqPiwmBTD+1FoN6MYsCh3kiD4JTdrijT5ZDTiasYh5j5BmJeEV2+KuzvisLZHxef
93Xh9z+J9my6re/swbelmYHugs7IWJDa5yAFng8mJPAHVuRnRBVVUiGcTlbS70/Hei8eBSiuroxQ
+HXkMGqGWKnadfvVsKSO7cFrS882WgoNfTPYt4Wx98bryUJlqf5WIqsbYLppGq/cGOrNBoYTnioz
Wb4qAb1ZCOT4zavE3N0B9wqEQR91qa+D/Tfl10KfQxRsX0yXVjnVl8DDy9RieQFq42N5UothRIl7
RnA0v5XOkBIFvUuk7vZbsG2pl4B8NrB+XZG+miVTixG9idQx2zKW8YxJ+M7z+yaDMJmwXVmAjdUV
I37DymkXJkiNMq1O7Zag182wYldYeZTn/9CQ3okx3vkC949jr6BzvzYbmJjOvtU/mdDGCPwzjh3n
LKUdRsij4doP1/RIkKtEsIBWG4WriYzbmZNwjpkNvTdMgSHhlgst+n5Dn9lTxVC060uWb1yhoSBw
OAiLJK8LCAhANBkx2l/+Wd/RvM0bSaYDGiTMp4NFVUSyYFMHQviQis1nOk75E3q7/KCm6tknvMT0
hU2rimV8w73np45QLbhYMSHAQO/jRI88tpQFl7f1c7S04NwL39aZbj7XF+gVDzLXxCGbpib2gapG
Y7qHs0l6DX7kAuC2+JM7SOCw+ScKB15h38zgxUKGJzOwn1wL0WEKfK9jEL6U1+40upucBKKuvRTU
KQP4NfgKjV/t7JzSzRkqQUm2JnBfUJB8XqvRe+NEmgvEUMZRiTEsmDOicLbO633cZ8gPemcEsjkZ
6X1Vmuoy/T64PpUo4jP8NFIatCihJCxPxRObBA7eeUWYjrNWjQNmPgJgzoHggd8/Om2Zu1k83XBe
4Oe1CUlsdhXBos4smG1WuX/U7sWeT9yZw4MupkS1gCcGWGFWGWG3z4i7sEVt6io1OtnCtS4DjAGe
m+L+ZtsRNin28fSSn743r2FD72OMgsTV1adl/N/qF8/RGpjPLMiPm7xCn3HGzVcLtqT++plwKnkh
G+G/MApWhktJb/AZbiuPIMcAEW9RuXdH2keX705A0bGblLHcJ+VGYPRm8Y6w/osnQxXeZI/4cN6N
QM+Y4Zohy+wlOFkvcPyNZXpnhJvKEHCTaeCoH+iv1oT7XNRyeLyICVyJHFaMd4m2aEQpf7+AlND9
kRYOomRlx2BQ8FLg/FXhsSHcEaSavOOX8ozrXHa++xT2XYFEYlRizCWXCGnz2DIr7R0H70wE4KnJ
7V9z3Ip/ZvU3yJcnwBihfFlB3OZsDC4iD3f6aTv++bMqspjrbaovFF1p5ilx3oXxmOb+E53YyrfS
NWNIsCakjyG8PqAAm3PBlcGjPPdaXZS/OL+Hs8TaRWNnd4GLSMcuRnj2rH5UZWxwIy/42cdfa3Fo
XIRoMIlSEAwI+1QEvB1AVSsATpJElCDcTUIfWpKyKHiNSMcT7KKmeOGGkxPqTKfx+9uBHvjPCTQs
oLcM25Ji50Iex08nwa0tA7GEh/snaV+L9bFvV0HY3LmSNOthKbFVKIs/xxP7PkOjEVxO+s2NXIbc
XMeG2C0LbNIrTayX+nXyCDLO5SA6+fhiEJKdqgU5uL0tRMWYuu5RQdI8FqfA6CM8s3TY/rVypx97
K0ZUSaDOzIqnTD9MFimH84AgmG5c0TT0AS0OtQaNokF+HlDf4s3viVromq1HVV1qhzbvRx1/DcSC
Es9HWM4d74Iru0QgBW2ToGFZRU0ooxqh5aYMsTpfPbdb+AiyrM4yDpu+9EQ867nAcTBcU3XcrcDY
AlbA87gQvi0JREhdzWus80N0NN0nvxVM0VITBdKcGSuMkiRVkX2eVDg3/qqPLWAKOVriwOw3+Y5W
OzCW2ieURYqVosHt9BTy5exOXTOO0+A5QCb7M1ZRKSExpbg2cwO31mYwCdK3i8uvw9VcWIZkGRbN
qTre/pgBF/wn/8aPPp4THzhI8tHCesv+iwXEqI+jiBO6cAq4RrY6HpAK7iE5DWtuRdy1u6yHaiSF
EeFzKlxezzlIF0Y2eZORr4YY5pXRvi2m8I6Buz90mHkzvvHTt/LatRWmfiN2UTZytKlhYNQUQ3CQ
ilawKl20JD8Ekr0zWklKVXKNCBaVN6hn+TbD5m4vyRF4MUlOAAP9yHiDRdPj08DxCOF8M07N1eTF
3jo0/ZhBTrlqjaOmidujJ8E0+AwowmMzVjY2efgbsLycBbTXERQ2fsM9JXYBrbinUgj4xLgg2TtO
c1LuIuogvtvokEqcpgS2ZFDB26a+0BFULYOCrlQ8fzfTR7LvdrLxFmzbap0KUAzcblyex9eLT/B3
owh/OKFwBLSaj9iSF1Dlcfwv1M4ipF4soiK9mDQaFu9K6QrV/jdwIsyiuaODdMAC9ZQj8mZKAEK9
D4kNyt+8OqvbA/bVgF9uAnii4QTJ1pDM2uJD7XojgTxoKbRPRW0V2wcR3nXA4ZUgfshLyPRx1CNH
OmQA2nuP45V413YfXf59WczqEwAttYuw6bWSlcXf9rtrw6nqzfJDn2Q/QSIu+3H9YH7tyCpxDSir
0CCAUtY/4vLIUP+aS24os4mJCLiFWa7Hydl0gjAOzXigM+1+iPX9g8m0NUXDtR2QJ8qIJOkBiP+w
I58ayQxRAEHlj8xZa4LBPL41QAA+j4wGdYmbLlv48NRIYOeCKkx6pMd9Cm7IFklnWo1fMKpnCbmc
LfYqwTHLDAiZPnVUZOEyt31Y2tLz2COGfsXtDiW2fqqKHnfgG8MrsnsbSThbmSAl0j9vX4JGPsc1
68bHQXymqyu7Jyxhw/84hqqoCVfmT00vh2uuMdKaN/IrJC2vzEh/GleMPo/sn1S28bb9WfYUXVDB
XTQri6UA9qbwLKRZQmiFKyTcauOPfUc8wnf7eXgHmcXkU+bxTcaAC052lwBpvhPqAr39lJHVfvxR
Q7+v+C5ndMFlnZFRGojWCZnHP68TZXfp43l3DqPPJQ94fvYw1lARI7wwgVgO3Z2DlsB/S1OwdyBM
EGPF/sfCz4JgE/EDEN0JGbn53oFoD733736F6ZBPiWoAnvnSaQISnlySJ7Mi/KMD813zF4EGEjW2
btTZGLVJ4F2JBiPuM6HhpyWFG9Ydrxiui3Rdc9WpBpVSmJZGO4qvasq39mEtq/aSa6OYipjVFxiz
Qhbpm1mo3OxoO1r2Ks4Yh7ooHZW8HdeKacIIob+WN3BqpewgK1LRGS3Q6tRl7lf2O90ULgicV1zT
i99PxV3Eqhlcy89eiuX6ii9rTlaiWxJ6U40pqv1uugBvdon/0USBxqWWHT1T3drFyQzR1qeif/O3
AUVc1xpKMkJxGfmSqLu33ZsEkEly6PcunrEFfpcs8bMnYAAqVcXha+nFjiD6PStRbrj4mblVSqtC
jb2B7DqD0YX90YgvNuAAx0Js2lGaplqTKKnUhSg3g2VOUgGnel+E6VjbsglqlUh6ESeA0zgF58b/
dxX8h4vr/KMmLNY4AnaQLlgehbAeMnymAUYc4DfLbthNR1f6Efa9QrIU8Ed3RFrFAGxRDbjBYypR
uhZ0iHByHloGw0kBSirEaGosdWbkQZKCT0FmhzDx//FrfnoiUAzworROxU+F02ojuLckm0XGOBX2
bb+yTJjBBmvCp2oC3IKUdKelSq5mHdYJvnkwxHQvgQoNi//t9tCrQYOYtUHyWpg3OigFqeG9ATwK
kYb2KB7KuCFzfBjUMZLyYoz/iJ6nLMZeAf4uH63maNBg3aHvruY2KYASIgpJMunV+YhlxSpszi+L
EG014t2OvkoXplQ8TWeKFiiBI4qcke957z6/xsty6ca0+OW8d5X65ao8F5ycJ6tpmENwzi/Ublk8
fahPRctDIHWRWJfnykA+lSo+V07KuaWqys9kn/0eeWVgQKhW2gv99Beu1JW0HAkYmXAZlIzQJAFG
AvCQX8UwWcczLeSY51PmaYxieHohw05GgTCZXI6prSINbEBBd8b961qwY16S3IANXgHnORfB6XKF
nAf/xmjg+uxSAInPvrq8g4zx4cVM97tvwRv3v1YdUkm9QVudWZLDJ07EezXUEZPO8CEZlXviSrJb
C+OX0txg8feG55yDb/5kwdfpNIeaRKmMx+EphQ/Z4Zoq+dm0dXl+vWUBBy09SymNfWNEVjlhYpSr
mqvoKk5xI1fiTcS4BW8OXz0/zu8nVplibLikE2DvYik6b12Vf0gQ4zawRikqNJWB1kdfPpTYkoJh
INfS/aaf69tl21RMo8uJp1VqI1tzyIgeyBEbxZp1nU1Awa+xdSWXnnIyPTKXSkq1TqtCRe1AhFSD
o8hV7Dbj/TDq3NlwjZEVg4pBPvQNv0HG6Db6+E9vmWoYAoWv3J6wWa9MnljTnVqhv7V8ZF+84FlO
n5y5tNQgvc7RyE79usq5kBR0BDbVF+8zN/B4lRknqo3hnHPYJHKPYIHPNUNITyRfDXEmS3n279nL
8kRQcPX7WIwgjV5BfVTECMFgE5Y/o4DBeQW+zIgvWVv6S5Rn8fRpQkMXcjXGEoehZtAbliONArj+
fs5T1U/E9RMP2Ooh7xWPtDvL8GhXNf+6Q+mf3/EA5hjDHSb5MRaNOXYhP6Kj8o5wu8Nxs6m25r/H
yw6DkcCmiWMQ2990TOqdo+p3G1xv7Zmzxote4SeLsanP52+C5hYfeYwirKL0pJgvzxr4yV1P93MI
jUWA9uLLAro3Ac3R+33E+Z6/NEw/Bdy8o/g1fh+p9LM+80VI5wWTTF07F5swV2YbS0FELD+SWxcg
AkzTtM0qnLGDYTWWRbMLE2wpyZGi0nxw4bO/PIaYCbqjZnETQLWb9oD0NRgiApEVDyOyDsBuN5kW
jdp/Mno+zbvUK8VdjAgGRownjqoSR9CI70Q24TigKZh95MpbB9oqCMl6jVmgGIPlTujLVkfxPJSa
lown3bJtCY6gXjuB2ozArfchNjTNlC5yh6gR57VCndAMAxjtXaY83O7t2W2err705aeuZChDu/ir
hYHzl4IM2cVY/6e4wkjvkSZAX/AobaNsOSpLz+Lgm3yr/MvGVe63Y0irjbGC84Vo18xvGm+M7njN
99aAwou4g4iOPSmTH3Kgk1L9jBJIRVemnfhLPyMSDWh0Je7hMAfU3XY2HTvzqa+OZ1W1cxPRILR5
SmdjojQY+ODHqSmCQBqAk2lY5FLkowYt1+GQIc8+dWxnuRb7pRKAlK3C9U5zSR3CWQddtrLhFchE
Os10/UqkKuEXjprPM7jHJ3+SHjd+HyDH+zbWnK8LLaA4HMYORBF8yRgxSNx1zmuks79L13dp2G8W
4IdBAauu6Li67+KA1eBpj4eRPTzbGA6LAFXujgYPocv/izNp5tnR/UQMW8MPZkOpp/iB0+Y3uPLA
OieRFH5+Tz2QKHKEOrsGtwatRb5sTsTaZV0DVkiJqYwSccl7R30ocxYPlu1kg9u082q+81RxKVWB
wGFLdODr8atH/liNAiyQ93BHc8hPxWytEUlWvh5Q/Gdo1CBdbbiWa1GmuIw1stJ6SgdKrObhQz2k
O1kiyg1j40U5F7MKWb1aBvLbOtkp0G8SXhyeyLqjlrCCcdFZRucak7xAAeA84mzpym/lN1PIN2Wx
5JVpXV0KEcmRAxwKDgk3LWp50cj8oB4tc7Bw3dSMTkncmXXv4lPBCeQH2qZhQYUS064hKbbKTeB9
+hHUgepwOJ4IlPvzhGrgZpmmjsMRKLC/n6kkF3kV3Rk9Bea25n/nUMjilQdC/R965ZeNel9m5HhA
9TtFgbBZ4UhaW9R5GR5I2TLW52hFZA5QqTBJjl2tZ85esLVYsoHUWN+gOU1YJgzbsb4I8ZUkDED0
ATZCvsY9al/6wVmTSZTXbiwVGVMJg6m9H32k91elLYCu9V3qrIR3fCR7JH9VbVlnU1Kwo53f3OXH
mRl5FMhaMOjPR0/cRWr0uZh2EtRABXJaL5EZI+cU0rZXeaghs5mDcrjkIsTfvKdeNDGjOloXXGEZ
/yosWYV4aXhkbcpR+Mw2+2fcFgBKo7DtI9Qt7zy/lC71S41JYg9pl5iyqs+0FMKHMliTuDz2HzZO
keq4meNB9Pr6iMfOhyF8Iooe/x/oiA1NWU9/uvKsgvg6C476brbGueHKE3SgLrLagPYFuuheXYNh
UN1u29A5Wb+PQ5FJh26XDRT0GRTFhXlbk23PwgannheYGUzNSL1nU422/Tki6qq482X7XFEjPA70
GLpxVIGPV39VfuedW4s4VdB156QBE4H8Pw0oj+qLFu+gaDgZFl9hv/dDa7UBmygZeXb7LlkeINfq
ft59ZWfvOhM80ihEc34QpQqSsZYU07yz2esct47EEUktGOarBnNSdYgACqDV6uIJYjfnjuUTDWN8
7QL9tPOhK18ws3menFiO97LFM8wj5O/IigzFH35h54+v3/CAHG/G4EiP1ujij2byiYEFP3FAwvd3
R8ZHsnIh5p7NaKjBKXMAzKWKCrR+3GOO5D7tbYhHKDdzq2lDYkcB9r4qdAbOvtu7LZq7LRfoNPAb
vrxPcGxTkRTwcK9FKjTs71Ser+RUAVK21gSm/zRVBTp8OEOjtNjRWUj9KDL3c3TiEbC0P8Ss8iSB
fm6pQDa6r5RCiw4LdRoXtOx688GguIB4YcwaF7/t/G6+MjmmiLVDUjszg9xawa0EGCLLNBEKASxu
Lo0vX9vbAdE5lO14r8giBON0D3yXb6f+Z0tpZ8xvdV8MMN8AJZvyKiK2fHLUrKqUjhoHWWG1Qo6B
TyCCoyhB4IT3q3JJ027309n9GqHOrabFsRd0d9ak5fdYmFkqY8pSMtf7jGo7P2sqW8tBsq/kLXXZ
HgMO5RPkQcESg/xV4P77zwScNG9bPCRzPJV8sdxkLRrLB7SIzXBoM11F5jFq2pYzt51c0hi1G+CV
CGSk00z1SFF3qXfd4gc3l7bdUFskcvtlJgVCfQymkwXfxWiX+vMLMDEzSoMcY5sIpzVl/ZiJr+jL
JxG3GOd8aZTBkgTWA1OPDO8N4F0rqrE5pAJjnP+2Xk9ahrWGz7lwa9NDB2kcom6ohEd2rJQdJdrF
MltTGQOHIIwSJ+roFTolSC7fFJ/o0815lWcUcNcdwO/DUkFjWJ8WS2rAYcBXelaoymxjsP/kWLKy
tU06UFik3qs6RYTfRff8HDnxLiuAXKAketaFjefaG77MkWPd5v5moSp0S78ETf5RotOrPm+SpseC
dkjBYv1iE3wUnnjT68tsyZ2itSHODq9X9zeAiTjVx79J0cn5lgPcWJMG9D00Hi0QBwNeMeWUItbN
lkaRpAqTpyL5VBzQJnG0KPOA+s9eRRSgdtt8xe9jIQtlQU6SHhRmxjUVqUz2sbmNvq+4id0Dgf1a
g7m+JE0yIA4vtvLQksWfPCDIhEF3+0UO1cySCvMr/ITEgjCx9dSFEMyl9krVgj/OFN2L3XqjvsmM
+By/GthbZNauVEmXkZicWInGdT9DO/ouLlMBJNGH4maM8Qd3JVnzs9JbdupqOgGTFju1gPhrKGl5
Kmg2qyAl62H2xCu/kJdsz51t96FM0oQ2r/a5MfmiEY4sVXpGzE2+QNUHfSIqdR/Y3KkfZworLh95
Hegz3j5o8k1nLOKv4Qp7b/bC7ypwrkJptEUR/oQDrjJ3ksLNIDt/wTw9Il6XGSS1cwY9FSfFbdTC
avk+2BPVxZoZ9J2XhyrfN3lzNRHe4Lz9nccVBxJtJ3FYFhun0APcgflJ0k2s9FLtgom8ZLHSsqIT
tR1ocU9olir5zTqw9L95AR+3p62UNget+Dy94tsFZXEkpKxz0fTJyXjL2fcfLUlWw4UgNEYTup/d
0xTuC6frNyFWc5JmDo3KDvYOHs1Hwvs6T1VgubcUvjxesyIY8/XPhERkZV5RyHzUp6ky87zggcA4
9i/70Gm00cBSMoQbVWGjF5AmrKpOMWGq7GPy/pZg4C5Hxf86rdvucWcfcMh279QrP0XEpdeCxUEk
ZlvWaKupy4ed5bvihLJf6MbtcWRMWt76MIT2BdtceSEfkPhfhg+ybw9kFNnuYMqQwAXdPo2xtvdz
9L+1zonUKLbMG9gKLaaFLhPan50eJo5chfyNvPbwpD3H6aq/AdPzDiTzAc/PeLMal2RGwNtvxSJz
/24ojXMAKMZbfyGTrSeceUssNlKmuZy/eD4ebJH7N4dMaRxykV91ctxxeF3ARJtxpg+PjZCOLlTX
34uEz6V/qU9aIkZUfrmJ2JepWksUZg8mOZ/MnDb67mQKNtKnBL+11GRCOVGeVD+lSDr5AIcD6LId
GsTglXXNDb68/Dp3sYumzhteBDIAbSvZFiMAfFjYr3n0fp0Z4TlJ7EdxCnxpGo4n3XKqwC7Z3pHj
1rJ1//QbA+u8fuWFyF3MwGCsPIbsNnjskBTQorrWe5+zvkyEm9yiVSJ8dxC92rckCnkwLm5VLPsC
zhT7/v60BleVGNQ5Wetg+qUuHh3vN4pQVp5qsIxdhCnphGUpfP6JKa4V83bIH/SPW6fF7UNACGDm
SHPnclAvAdzDlfd3APosoPHJWKRAkBmAu1baIV3Rn4cyrex4D2fk2ekhqzQQ2JX6hBOQ+YSAHYIg
oQHm9nDkVL+amKPq96FatjNbkWMscU2mNatkscAp8ybQ17tAU0RUCYier1KwBICNKJRrqb4T7Xzx
wrw92kqpncgmzl1jdN0Nln2NHfi/TfxXta8TxER4ozlyndPilm/am3QuzDncznTdSF7DEPZZGSru
UYtDEL8gVPktxDYg6s8lL4M2kiNZDmnrncHqmAavojgrtfGyklCpmYu7iNBCRHE3ulpza7BmtzQk
AwegsctkT7JBBd4aYFEABep1AhGBwSiaPafNIj6BNROUOvpXSF48K8U9GVBKHrZOGdaROXZvB/Bt
Qf2fdTP6ti9HSme67FpBvznlYnQi6GwDOwfi/4ul4MEr/iYCKDyk18EFgTk7joCuKLf0SX5+58mx
sPKi10zaie1UUm8GeCTths4qTWIwQpgLJ/SqNXOuViNaw+3nYZ9B57XqrhpCrVcn0pYrW7jIGMFQ
QnTW+WYQT7Tw49rVoL7UydWx36/tt2O6eB2VD1jxYBrOzbdYnSjvdWvkjYYPHs3rwmw1Qt/P2ChW
sNwLE9Efqcq/UaFcSn8iMBk9ANDj4PFA8QJlKyF9hpKzaHZb1HIJyLxJXG8aOOk/yQCofHlmCHQN
MSLbeUQuAAxTL7VNColApzsVsmF0gxlPfkyLvicF3ru3WG5Hc3PTzkgKBVx+b9RltnZZ2vx/SfXJ
RQB7Re2oTJLCEBCfn0WjxYxM/4zclxDOlosTugZ0M7P8iCMHeiyjrqZ0VZS3QxBFvP8JWWQS7SBW
4o2jtdtBmGOkMFQ/9imKr2VMAZVIbTMrGjsREEuJ6rd+10Yw3u8R1zA9EMfT7eSls3oh3Jp64O0S
IPdLJW2K2ES5yB08njGyI3X3HSkmpP5Dc2qQ6KC0I7NWb5ot0P02N/37OkxLP7jkcB6Rl6R7EAHT
qNGwNBVq4J7QvwaPdw75HauCIaqaI/qi0gwTiikPk6L92zIoyDcE5l/WAEdvJ4Isk1leXSzWPC/o
YJvC9P1odPxZgkpQXDrnX9GQ0y2fWvcEP4dcWdt8N/CJw12ptpbg3q85kAbL6lEhLNyjYu7OSnyf
4SNWPDkNJM6htc8J87yrQ2U1UJsY5QQp32pjxab/anlcb2JLFczDwDE/SEQTwov9x2MvQp6AUTJR
aGpenIpvMgVQlfmC3BZ+7S4Zfmsnx65CGyxegsOfagjcFn//Motc/S8zP2GYfLtK79Mykre+RyZA
oT5lkmV7/kzsx+2EBA/OJNmLmRT7bD6z+QNI69udksJVik7QS4j+PSPEZrV68rduioDx5lKIuUlw
ntzGH3UgRtZaWw/n/CA10BpcbFifwe48IPlIo5IQPJazwD5r5UaRj6doS7MfiBEuUUPOMi3FTN/2
enf9aadjZsk3QjOdLHJ8ceGvHU82cv6DDcdikCTDEZnsENYTTguE6lfatXsVcBwvDimoydz2uIV9
0j1DOjtzI+Aro2koyungEbLlORo6IRmVkn+C7ob+mf87j+ZYABLcbmqXUgXnpjr92VswsSmT3xmf
gWYvMQE7HB0DpDRgTPHvMy742gb/XZHlqsDv0Atip+9RUEG7928zH8EWUmkNb1O0m1heVFzuePl+
A8cph1FCgLZwoT6smgZLK/klD6RhkLhZY9YBPPRfj/R83mmU+Ze14PpU2so/TarEhAcnNBXPn5q7
v0ADDDrZBmmHGQdNy3jRnBh5b/GsBOSz3OT3ZDgMqzMrxW9GRBpBbiuAXejfSB6sFcjjIlZzGb20
b0a7hc6x/F2hpRJdJUdJyT/vvWVwgzC9CZIOcvAVIIhz+bJzLS/egvzhSG5FYVwRdvmqp1HF1CsE
NtEf476aSCbvZ2iJsv1uAGpZBbXhpjBVZTfcu99pfnAH0i/hEyDsQP657i+4UWm7q8SPtIRekDsY
Sd/2cIi8XFVNHYvUnZdE5tvvgaA0IrZF+bkD+9ilzHYaOtxdfDIrXCYXknygGKZIiPTad48JdS+5
Wv00rYwkRks/HJKyurbqzBh3LaQElJF8LhxhORXHeImn4c2AXRQgbvPduJfUbH9SwSy4SeI7rhe0
P9YXzHIjtbq8ZczKHbmJGHwj8fdguUtQKEb8r2XPRbJJFrZFYYGxRKxcIoK/k2Bbx9kXBjU6PVCy
pVjeqUNfLzCXFuH7QZLqOe1rOh8J9w8iXwGYeDgiFm+XYuHQSluKHVSVXasV+RygOzNCq4AK/8Rp
DGJ1u37DuPfyOQSvwHSNkFFpdKEc9LaIuzPfxBgKXfOp6Zv/zeZ68SNVZ1u4Oj08LXPJ0+Q5/0/x
iq5ngh287juUiC4R+1/L/YNF3ZDO+pgWq6DCG7Xrb/1JZS2G0y34b6+MrlFsOjzH20iRHOELKynZ
Q2ohMqToIiwwc3D3BVO6UHAzVWYaGgFKotgmG2St1xyspsbZNAJ625DTUMxxCgha6WzAu1vxfiGU
0ZWVrIyPsB4Av9hrv8rzFs2360haWJgmi1Ml6eHC7toVo0cQuJJw7RjCRR9W1o3nhjQZZ3tb50eC
lrPkFxG7A/mu2kctjCs+X3GrGpMSWz+LXeNLyslDTotn+dTPFeSAx5Q0TZzb+g3R6gUvr9YsP4Sm
boNxyV/dUXp8lt3qkKy5EAlytCid9GLTJTiT6MNcBgdEadd4O90XqEIw5Xl8rMaHkB8bxoDvI614
HJdENcj1VepLMHrWyy8FYbrA9EJ0aB23RIFiH6HeMc7FDn131oOYsNIogEJ6jQ9FacX2uPLo44Tp
YJ1rufRSIegX54609mWanaMe30gjoZcWFe4+eHn7uYpBPqW33UG2QpF0lMdmEMfKDd2hBQnDfYo8
jjx2RplFwZ+GR8zxq7odc83PE5igArpEdEyXhAIQ1wf88F/wnVEM8XD6IF8BHHaxQp5fr11dhAJF
3FpfTGIHwO1VW/cMbuGlx/99rJH9hbgRVe13/p6paN1Alq3gtMU7g7MyezgPeck73zteednpzJDl
D0p4SOBrhhODOIAjElF0dtFUtJDelK+C7Ojn4BVZFF/1ZeJyHX4Iccn82dKfTblgCP902ipDjFjq
3/ATr+SFjtGy+b+ajrIXszcF3LybHhKh2UyOUvreCcSxaRAuUHnC80UHvlOiCEouOw/zlD7ne2rf
JWpx3dEkUGmvP8L4qsfTF6x8D36nOm/WGORl7MxaJ1ZecdKHusdczCpsyP4fYxpb3x6vb4Uu4j6X
tEHxY3BKRXfSI6sZ5RmpRw03xK981YA+S2XJn+F8dyZyQYXB7X0G2qC4+S0gn2F12ZdvaSc66cet
HJbdQ2qKPa1Cy9auSoBJcG+MIw9s8C8Z59NECxVeOJZD8nN3XF8zzCdhzmJ7ZJ20wKLRiRn99zlU
rQB0vFrWMPHxXPbc/lbev4PFT+MW1DxPuZBaQ5dtSzKz2bb6vOR0WwZwKEj6bGoFO4N0IfRcYGdL
73MVoQ9CcukAeoe3Br6mqVAFflP3nJtgi8aq7e6wBLljm0RkvY5Y4/SxB3se5mwuDksygI9gdrfs
C5l4MqnTfMl+Uiaru8XP82bd+ftq2ypsZQxHUL8inlwH/X1S2DVOT4LiOJ0lZQW+Xa6JKUzrgp+r
Pc+WaLnlxhA7cafQdSgqph/mYgMpsi5hn9l+w6hFHmRdnOFkvBxExXfTMq5mgcnk+Hl+1rEXSg0P
MvHkSwFsGKKlvTDUajWlW9s09G593q6lMTcR7a4wdFd/X28uw9cxQiIAHjI/vCieD9lY7cH0Z9G3
9ZiRz46ffEEVMbkA85gjCYZYeF+iygpoPSKMy32nDWNSVlspgmP/BvKJm+WqTrs9wXnlrC06h/GV
j8SzVMAZXoI0KtmF/yZhdH2fSB3APspxi+GiMRLMTmz2V51iiQF288BtF4mGHeiq1EMDLrTSuLaw
4qKw7c/BPMtdscS8JBzojPWU1YnsV3jvkbXh9OmzGRM+6OzUMGz0+tFJi22cAeYeY3OW4RIiVuYF
S9ODuqdzM6pP87nXU3tSXQEtzciNvax6giex0zQQG16oiKzQy1rG37w3CoQKZqnUCgrx63E/0jgu
PsIu6ZWXLVe9hBQAImHr6hJtt+6x/jJgpr0YpsiThJJjI8TnhNVRKb6fZCtgA8RjiQ7GTdLoqFax
KEYc/365T7+99b7pY1fuVprGA9OaV8Xvr3ZEy57xZmVMaywM0at2zhccVxE5D+yZKPcLnEYB5FQH
SuBYbJ2ezghFEMdO5H+g1B5ztf3Mw6cYqPSQ8/B8p7dVy+27YChAz6T7cyMQpwOjeYKaUiF1g7B9
ybZqNmoHjLXW/3LhuM/ME4pM6s7f8TeO7u/7RhSxGZvfZ9WuXv5UBva2o9IPbhcf8b0SQZOJZool
4D+9lutYycH9586uQNz2AsDkyc3YvhrbMQxttEAsDWgNIzhtKG1xFg4279qKTvOgHw0LvXkE0T0S
sAubpDAVBr9Cr0z1RNjV/zGBo1y2EBqDMNFL0/UbMEQvixsu0PO9tQFt/7J9IN+Nm4PODCQ3XaQf
V3pcQwe+WaU3sSx9aDbTVXnCZVOO4G6UZXmKd5tQEQtuYwTuTcp6YoOkPYN03/VonPh7g3+4I8CF
jLDDIVlWDeiHcy+49QPMttgQv+J8ltfQ96ruPRvX+2atLfORC4geteET2Kh4t22DHHVYLETC5YyF
827vlEUSqemnY/CgaANTbroE2fEZDFqY9+1IXFdqyFtmlR995VyKXEjCd3Oru2y5ZnFKh1HHUYUZ
9+HavNa3CkHqHXJR5ix5izGKIke5OqCLgGpXJ+wnV2gDllFoJGIw08kuo5zGbAp3MAKrdmZhZhw+
oPh1s62cDHlEZK6vW7iXn2qj9c+W3IR4tbfha3FhF5Vdj24G+hX6nwfB2T+e3cfPfDlvaVBy9TQD
4bQKi3+gm9oieoKjKvqIuxFPvfGdRPhKi+x938yAR27ZgSnDUItgvYBYWjZ7bLsKU49PbfJ289c3
hU4dReIxZdPjvapx5+vBNk6NgQj28w2kKy2xCGGr1ZFesQhezR+PY5phS0w+XD1BjgQut/EtHOYx
WJJu4K/J+1b3KOu3N8Ax+ea9OVlpgvlfaQjapLtedYn5/xL545Fp2aIMz+JCN1mAo6+8e4U/nOU3
orJ+CHCSfI/FVH/cnzMDQPIQPHr2sQUz/mO26KCqsRfsDRP+cEAXxe5bq6vubVkVRVX1qUDpBpwx
z11dD0Txa+6Uhol3fqFawnLo/xNS3ewA1qdWPqPnTCXrgacmIZr6vRj5LksFs5U5GN+FjUEFCz3T
NijSHrPCmaUIBdAtcjbmPSVuNdNZ21yBn/Yr9dGzyKidsagwoJWWD9HQVJtjGw73yExF0XmsmS2i
Z7uU4gwT+xolCyQv1Y9fzMxEZ2HCds+FivO652xCSOhgAti2VXAcHtF6BjIbu6ZXaQsVLH+1hXRi
f3x8rJ+pqDE89+XxHt7y3yvPwhz3s8UDHVb0C6Lhm4al3MifU1aM8BTkhTxCEaCmv9MZ6g6z5BOp
67v5x1TE7GMd+d+uDl1o4czROqfj3A3pUsfv+mcsOsXOdTaDOAUJt7PgUysl4wTmFeVWn6XKb1TZ
+fInWtw33aW4W7UeH0IHWbxi6suD019M3EOYXpVrKvN9ydLoXsBMPQhJx3OImNl9FJXfGJNV71sy
i/QXADLjyd7u4UV2qN4e5I6ZOZbraVGsL1Q3ZSAHUw01hvfYBxV2c400xglHD8uw8P99+ONOLJpW
afV9f/4qvnqFHCImniw/4BQHtlS4B5x6zTiiLH6yovWRM+HcBSJJVp5i4A9SgrLQ/ETy7zfiAjO/
jrskDnnr2BZ0RS4RzIP/w5S4btU/YDnfJDoNliK8E/gVtXsF/YZ8tMvLhZQqORigb0aPWSLC10UL
R7qJM8GiNNiWPiL03PnA/IGGHJI+xXPUw4ToT83qdbQqOn1/Gj9TMdZg6iriAiHFt/mOSpyGPby8
cQF6Q0JgweAUpQ6SkechTaMawQrwKGnv43rBb0KI8lDs9gBH8Jd+ZJQWqpgEBjP0MYR7TPAapq6R
sm6YSYO8lBtUkWhpsvbBXS6Em5f2HC9JD8ljuHFum6XEqhQMMbjRJTSKlMmd5yLeI0XLg8vlQoE0
1pUiDCUXjJ149dKvApsFJXGntu4/9RE3DCJqC5CyWq1ieNaBnsg74fnFND18GyaE57fUow0mHhsc
u0KnOcosrAhzFqNAE7kFtsFFXF755y/W5/dFsr96RJft/1sLqgiix6d7ls+p4OL6A88k+tzsiA1f
UVTtHVQZ7PSKTo5p/l1feAqzX0JCWaHVxVT1iXLZtBowxmHJDFNMZZe+5jWKp260FE1NIwLyczXZ
Fsw7SolSaf+Xql8omnFt1GQyslEumY3pfeVt9S5VDpy2jI9l21NDOh0vujDkRUjhtsNuU//h5QGb
dgf14bgg4yfxihpUz0puf+CNtChZOK6p6eP8cbtgLNrqQxZuo1KhEjHazXpIXUmlGGuvSWGr9T2z
m0DD+aoweu3PZ1HZLyHoxUNhYnV96auOmDrPgy99wkjV+/OXN9BKjakbJzgIUYtYRhoHyHrVJdaN
NOQHr5L/JFahOxGZakZT4AUiRn52SZnehcBt/NA5uyuh8T9p16jH5qcGJAyl1gAnYywNj9+8wCT+
N+nQlwJB4gHd7OBtZC9IEXmCYPRhYJC5/wffavZtL5WAI8NCkKUL1JeVjeQblLHJsCafmLKOB+qg
jtiYYVzX6T3iavH8dByLSuTok7dqWjhnhZtJxMY1Y0FDGbWf8mSpX7qsLM2riGvvRVbiyMoXX4X6
aH966Jly5SJtZ7iQMYLVitR9hS923TT5kAbfmvAE75U0MQIx500SB+0WInifF/JHTe9RABmdyDFM
1qK9nWk9RxG7vb//ZgRMh2L+z9FxDY07RxFGUqWMQLIQeC7+Zm/U0C+3fX0oqsY+ZVFQ8HRD+cih
+G2B+t5GnjN5qMOOcFfxOId8klbqyVuvA4QqxETpAHbytxwhk77gt2l7XqPaUyqmM2GjPJy+esE5
j6qEeaI1YHIWbPx9ZrkYrFI2FiXaKv3JdvBaSf0x2y5zQyyNmcBRevMo0oeFY0RfyaAW98dsSUcn
8dtdzVdopNnh6afu/rIwK2T6+ywgY5mYnsTtVtC8BlmROKPjX291BCSXN/AmONTTSxqwihG0DGUp
Z5bvE5u5hXcOnmX+in5KtJ73IabveeZhYnJuOG1T4P0m/v8xopAcnIDQGpJH2kGxX43hWQFXqgNd
0XPOUvgIWrYSqGUeVEj11sARlZvXrjNkXJ8w/l7RKAldXob2kJGLQ2c/W7Zswx35qPaPreKdCHt7
PUEtQWwJBJZRalMWUC7fkaoezl2dXRNatgpnBYWftUi5xXbMs948xg/yRlPQPGJc0BDPZ3QR1Cuu
2fK3kLDmr2GktFH8vZucJlCxdbvo0Z/1jTSgbkdQI3M5fVQs14bl4Xe+a+2FFJfdY/qZOvgBoC6x
Vls5pu7mN3EfzabqAJNttlWPN+eOCcoVxVCSyWAWn1rjBNWlyRgJcUbYzdxBnUHz6a2WULGh/2PU
iN3Nx8zGNbAiMgK8AUSeI381Mxloc9blgsY29ljy8mLsNAC+xokWbj9Z2U05kaI7Z6X4WGb9Fkyj
d0dzYM+wfdN5rBwCZRwbN1UvJtdG9FMlUQZ/QSjOzqvENLf0DPtmZMXnOCDcuSQWDopc4mmDN011
NKz4QQJHFPswb/hniUlUQvINDQizAp9esA/cnX3F86gH3EGyy/DHp+9LvNYfo2wZib8shRREMtxd
4yxMg1xDR55abnPZdCx1ZT1deCqpSIzoI4xpGDggZJ/uZ+sjwl+4uVTn++dBGZ2y9in/13y6AK7v
NMQJfZUzllSvELg4xbydQg9EX/NCTkRG4aFw8UVL/smmJ4Iv/9jRUV2xIvbPgwEN4VUf+ZjnqeLp
gk5/ix7OilkB7gzMj+3U5xnpDjCpYIxaSUPU/91U3lzWEiBmEXNUwj1xvE7oOQMBVuthILAJmq9x
BDkl9v6awzu4W0I5Pt1OyaKIDaEsbtMr4JDc3bB7mfJo/POoF9Yt90g+10bovDxqqi6JKrGHrj+S
HrNQ6DDHD/Rrz9+MCXSDRy871Mvs8LAg8wZ8CosSRf/eSEPOf2ubMvFv7u5TQyDB7JODEVgKlxwE
TETa0VnQ8oG1Irg6g7yEYGQmE3TpdfaT6BS5AjhTmlbmofSKBKNdrF3thXQBnjTzx2GlHLI3GtnD
odMJbi7A5x9c9mYsXbJl23MtlMnTZrtDRUuT6gixCbWznEykhVDNs1mVLTWRl7zmeiixi9OGd2Vn
gLzcfAGJsC6EqK0fv0Ivsq6K/FD+4ht3GnwYfJi0ELFKk7N7JlNT+QZ4pGCB/ZgtFqAVRy5ZsXAP
E8+xLIUIJTwA/vdKpBKtYTfhuu4a2u0eMKvZCMSZZdFJqfvjl4xognh6VGS9LKXTsx7sN/XBPy3T
/GMPSr9aB5v/dHlUV0bwqf4AgeV7Vfm7KhMnyc+ilzTrZo2T+TqaSkNGITKihj7TMjXprt9yH7n9
2cNpMhDydy9lcx/nrj4RpXbfWWizWngt+EjHGhHlnlGFF0+Tpz0T4AsKQK+YtlyAF/9xZX1TB4wX
85lGNo+05i8ghKpzXZqWm/5NAanoZhhTld/ds7sUaRpSWT75d0ywOh/2ReG/52Im77EMjkGC5nK7
KB+MqGJPx0fAqCiM2irOmU37Zr3nwyAQvakNr6uxUaQ1XMLUKkhTb4x3Uvc6DK/r+d68cJclZq3t
rMFCubD465PYMAy0FGNqBM2MXQ6tkXXI1avna76BmELU7Ay0Ty7wBYLWiO0ToIwVdUCKLHxBHUfD
5oyfIPQfDN52+vzi7XSDMIIe2do6Uu/Ijal7taM/e2HZg+a4kfqEA0vRPGgdckVtNNRoFjSgGd5i
/t8UsQAO9+fDMzvesBeS5zDEbfjRLHv+R9oQG0clUwcD+IrSciqzrkGQTNvbvRl3BRP1cdcgr9co
JHKD302OnK6YXqAJPSoxajbdRDyXoYlMw0AAPqY7iZK8qRpQghUQeaFcC13oHoJtBm0vjFEBXUON
WAXiGzPcsbYNBcXN70RxjX0jyox385WCqKSbqJ0OlXuWub1NRxd2FK+cygjA6ED3qSDuSbcWSyRQ
mWweeyPyEf5Zgei4LqPfL66kYJDQ5hRVBes/Zwa0WvTqGUBKhlaRW+E/gLFaGjmcucw5rb5QS0Ru
iDg94BGeGIZ+1AuVOc+EgKFLLUuVRdFBiImDL+WFzg4pIZepNWeZnLMNUn3UYij/cO0fyJ673Mpy
tPttBGccPZtppZ25GLyoagKmvdk1mYsi+hgxdQ+4zLXo2Dkrhxlcqyn549ovwnJzDcKH1Vkgd+Q3
Wrm4s31N/2pRiROaAdIQm3cwvFyAnho2hAbwaWfFHzHS1wdj1Ej9Cvsmn/pigtuZnXDQj3R3gxgq
t+jdBaeKHj0e+A3RJNQWua74iji/W15L8XguqqCw7KKq/zHAPfxUZapL8hgeECym6pE5uU4oKOMU
KzEaNDrpEZFzPeI42EvbuGmnQzOUzGGxyofPimfwmFzaM8SfJ9cGX5ghy+IzqjS9QEysy3bxVdlm
3iuoqDlOFdBEQ0Z/wfp7DDipXcfy1RWzBxQrhJ2vsFrWvbAILIhNeJ42WC8156rpzd7lE/dinGcd
EaLv/2cTe2Z9bcebAYkQpjLNRN7Um/443CgfKDQdTzA/G43Sc+eSB8hq52wSYuQE7Ke7FcRI0Jtp
DzvYjOObYL3ryKw5jhIKYaqYFHTovOlUZd1O/gZdD73HbsSVE+NgZuAA34XJTYIX37c16ZwQ1+hm
ePTbTKC1XT867JzQhaWiB5VkwyzjNEI5zi/mXnqJTjDMJpr9sY/BSXZw8XAtNcIotxGamFwPXnbK
savo739+RamlfuW/5TVTMRF2k4C3YQA/33giY4eXKhjIBcZrOMv8LJvGlRLDpZkzX4cw6PBeegxu
btC7658yhpstjyQOokbxUAKBouesk1wFVLtfYvKefvz+1sbFwqaVAUsRLIiqJS45BA/Vve9vPg1U
+L35gKg1jpVZNPkESkrmugjd7uurW2DeT0P4tF8/49ZrUOEi6q9LTB2hhbOuhZCpMsZvCLYHLHYX
ZIwaopegTGchK1gIJpPuDTuehL9aXj16gPx+BeJItSV6wIzShwabf8IQpJrDFmG5/U0YHoKpOkTZ
WMxXpEflhFRMOv8Fhk7tpOHwfDXfE1ID8TAwicjG7U4yoOyuqaEDPeh60nD9StA4y2D7JUEYPz0v
NRpbpqVtb3XG1ic/axUm1s7oEr89OMhQa3aM0uF9yDmYOzmXYrjXbXjbFGaL32tWibLhSCQQ9Hl+
tcFX1vXIc1oXK04u9YNoqYdFUmO9V0Xk90UthwRrXYzvrWAgrg7mKsmn7K9iS76ZpczzmyMD9FcO
JiKYTCB8oMiDAYIlTvZAIz4RnOwN8UkpnnPL0ZJu5MsgxSmxyP1aL2a8kFoCjWbLgpc/9zQe6Iu1
koPlCfh5AtOidyT31J1AZwl+jvCVj1pUr2L9FzZBSsLmwgWpfUZAWA2qmkPCi1GemW5400V1N1Fb
Tob/Pu/+OgdhPF8pklkIVdqaQrgiMqp6Kcuf8n8vihe2VX7HVOb5/RLrecR5tyszx9dq7m5Nsp2R
2XMYI/T/41mg9hfGgyFe2tdx9M8NnWXBHCzaQjXh20vG65x6qUUaW58wLKFPxK8gGGSBL0fH2pGv
QziHtqabW7Z9OEmb9DTk0LPEFAa9HlCT4nJn+pVw+A5FMno44FecKHOvNNj8K7KMQ41j7lvCc9+R
MPMyU4Zfw+paURGgARtKhGu8l1wDmxvoHtU3q7dyu64W1vtISLKY6r9ERVw4RBnHlhRGILS35rRP
jYkCRZ6RMNdMeBXPv4Jm+pRUE00drGK1yakDv8TWs0qveI89JCIBs6k/Y0kpG8WmkHNrlwgIpoRA
fea+Pls5aHQZ2QA4dQws5/lMoL373wJpyNcg+aqXBl+FIGw7yYbPz4JtYJVLOE0/FzEjKsbsURrW
tCHQrIGfKQI9962qvmaTwRMalnVNV7r1QbxtOD1jn3pzLLclgxWCibXELXbfoSFZ4XFxFhhpF/NC
3jvsWSiMIBkimXa5rDxTQkumZXgXMRlwTaNMFp3VkGTW4bRVijBsH0CYm8K6p+0qyMU8RddNQFBP
5V1n6zS6M0S2bvNUUEi7ih+ng+/I3io85AA23kZ99sk173OU2ZTzbBhL8DenBs7t0hYOaBM6dcY0
cnA1eothKWeqTqqjFeTm9xyf/ITyBaZG7/XbDqwcxcyLDqZ5BcDywV+7mFfgpYRF4C36NszdjxqT
OpyFahT1+GKm1uTXZeU2ebM+e59aT71CbF2ydJ8JJo0TflXDZQpUi2rJs8AsMIKKRsripp8vMXRe
dA/tf1n0Sd4KrG2uXx9YkJm0cSTyHILDQHgdDaLwQNs8UVzrR4JBQl6Lmo3JB4Qs28JNdANQQWUb
LFpFHDGKjffyZ0hBI1zmYkeKPyKaXgpGEicmwSB8U5wJyiRsVzl0eVN1DpNY/QJmw+6QlNSJE0tj
fNaHnzQ9aX5bOYQ4CZPIa+x90N1UtAPNklp98h1GKEPLj/qryzaiydxja271b2o3qe4k6SnHD/Mt
X0IIrQd1e6CsuJtnakjdmKyDggwBJ/hrx9xoqyTxtTlYXeHgPNLEX6g2s9LmnZOH5fRwk+P0xyAo
eq9kzQeP+rE9K4/+PdCunH3E9MOS69GcWGlDYzrHQWplOFt5bzNVcOnl8u/FnqMJdgud/YZ6LDEi
sC1sM5P8UZK5mJWuvPRycFV2RlqRZh62EO/LryREyXA3CFPO37Tubqt14i9JHe2P9//ckzlljmBv
yDe3EZpHwwgvKiWzxoA9btjl3MKr3LYRrAkh59dX59GV8f+9X/OHOkVQnzLrWhZXDOnB1ILDjIHH
dxx2tVf5i/ecoZ5t3xqe8BeHZiioFqwRo72TrvcttqPOosbKBWLlYcJq1iuuPnpaq/6jXJl0dvgx
mpSM8MLV8atFw9TjY7kM5hjcMI05bFpWAo0QujZmtgBqlVtO6pkVodkQCgWVpdSbujMJ6TlDPxKQ
Ov7/r4dSQ5YE0013x/Te1fvmzK2uXx0xO/URO2yUTWu38mboa8K3tSoL7Locb2bMc+dCGJ9uAWf5
XT/IiXoC35MzjQHG7pGAocza2fijIK2439m0yB6FdW/gCeCi2qu3oHIciHL0PiYWogRTuQJtYq8Z
AL55gDa7uSnH/4/oJITNVdhPHrDzLHOypQgu5NdQa8pUHI4Oy55VJfOpEzEs0tfyEuc/d7pEuYvN
NSRBHt5zW3k53rqS+XqtJPw5NBU3/FS+xnvjXQUIpH3LFXvlSpwIA6eEM2Rvzm+y4EZr9W9t+3Yf
f9QP7eJwkN/xX1zh5pnS3+GXkLHDTIC/dfXlsPehnIdtCpy538XWyXASEXHKhCzPDccabe6ENTjQ
d5qntoKzgLZfzb6r5LmP3uIhEyPilk7dH2AFantY97s61KLSlqdtqy0Sot8J5o6EJM3e7LlQ7azv
UU3yYE7rzFk4KELeZeCszqAlzZCzF3kbLpDZVFkSM2JghGsUaQ0+/zrE6kC1LZwMgXxHQ3fAVnMn
kVkP3l6AbV3BKHx4MuB0OnZOB4RysCsz8y1du4uNQPAACQzyrlnNK/U5nPIs2/gP/DBq6vHFzc7t
Kk2c1VP1qcjaJaA2TCHi1S2zUKKNkbeHRlkv/8OcVjqo7xsYtE1SC2N5au79QkxFjacL4b9oBtST
KIy2GlSrb2PKLkOLVjxNqsXZgodwhZfsYnsP9M5kTZ79DogPh95XLEjU52EZLP6GINH7Z2q0uTyU
/Nj6xwotQuSxR1hlYS4qVLANesSOweCIhnzyhkwyaxFaphFch9GOQ5qyyydLKnHVvQrBR4ydkWWC
sMcC8BimAx034pRdwYUvsGHMR917ZkPS7ra2eZJEJKrwDY56yzHxKu/qnC4cseNkTP/4NCUE8/jC
JVq6b3VQupdSqmPytrGo+R381z3aszKqgQXGGWp6vnyyzEuU68/P97D0Ek6dtabLu1K5lgzc5Zk0
90IgyCvG1z/D0muqx5/1HA52Biph/MKiYi7R7ABbh/2EQWG3zHR1w9r76S0JUmXsr/Xn0UPhGL1p
34hK7vC/ldcGjt1VEwkRjAaEplLxD2Hg9TbcfQ2A2O8LlZtknnsxNzOvPxlqUi0q/va5PDQJufF2
hcEjJabm015mVSlVj8S373ddanvSl+ICRADXfntPGPwl+drqktRibIqh2zqkzl1yyDUci9BVEuxX
Rpt5C8etK6vbzX7x1h/lPF43DwWPXlykJAbl7Ps6YKw9Dph7wC/b82n7kqCPXZe5L/BQ3vKZcMDj
j9wNh+A9AWpZNvTUKX7lDKzCvOFPZTwB/T8hPExTX98ugpfJMWq9u62HtKt21nlRU3aSFVLe6+0G
Ubpc4WFbdeVQL3zTFK6TfiyQwOY8IDkcIgjwsLSx26mFtlBr3FnJ0nfWZHJlbC55e9D4VSilh+Vh
AED13GDgJhlvyX40zRsrFtJLlD3JGDwPGZVppXgWToKh1uB9I7AdSKV914iKmRtWyDtaII5Frqo/
Xitf0PpaJNe8TNYrQXZvvD5BElwvI4IpvugF6p2kASnNHUeSAb2//wFg7ebrHyZnjVLO9i6wwunM
ZvlAWbfnUVu307NFYpOlMXslH9ZHMC1SoEu9rcx+d2USgS1NmMGLEpB/Zrsxb0IXiQ/DmAhiFtP6
xHKZXzAcz3Cg1tsal5jkk+WIkd/Y+9ymQIi46+UQD4VNr9uvMpB3t4kLreuPs252Az4Yyo4a6Stc
3l4I4x0Z/3YZQFnWaa7jO7lPwnlYP2YW5mXxXW9g9YWyoFJwuhLvtGtTgdkeMoCs2kNFvLfJjdFP
LwK9FYizBMagaOW9XgtuQnrDsfTYvJducEybt58ETXTedzdWZMhF4vk1myRtCf5nVH4NjYzkFz1c
bqFb2GkFHlis3cABk7CF98s9EQ1Tf8DhZ+4eDutcA0TbKBxCOPXaUHyuA195EwtBhxikZsv7cAxf
lGGnMrlEcSowlrc4UNUmr6nkTNXTVgRRmIRyZnFZ4mpyM0anRiw+pQ/W/FDWZLPWB+joWM1MbqeY
rpbMG4w8JrLHyl0KmwxE3mEv/n++JOzs2xhuNDWo59nclRlsj+qv+ZKgRyL4XYthvogDxCwRcqyB
fVlFTiCtBOjc/VHAE8yO/a6MwR8kSL23Bil7VjVRkBrsg6ECQa3Gks8//Ejuds5MIW0+RBkSd4cY
kg0/WGCYdkDlnMKWrO+nldWkIf+sfofJiCYVPWTlNMcIGXjJOuAfk0JtuwBGtMYopcC0loSvu3dC
n1ya6UG3ZZzAS7AbP/o6k9Uk1uaPMipOW3eSRfUeAvXkE35Bt3IMoMeKgCVBWFA1KQUDYYDWOHNI
HtHetZSAJMKjjW+U5opEmqD1iC4P6JGxBDJw9pgXx+NHWw/C5yr6sWDOv45xkpI6itJUh01E4FnH
CPHG7Cwrauz0pG6JvOH/kRuvPwYXciyAC134pjXCmRRRLYaRa+/mTacqVY9cMRbhxH+fjz2RBz/K
hyf2yDukWUvREn1n0O2+6Tlir1FEao+3ih08oaWla6d3usTID2kj35mQBc2lCQrJruJIYQlzwlAK
tZxHoUCVZjFsLCGOCe7EDkMzO+14A2Lj/wOESb0NIIqUOWoWjM5GXHsYfsTsPihuDsHlMAikgxFU
OEqbU5ZPBkoc+rMna1ugydk8TA0awhMeJH2YrlUZoXPf4vZKWUKfyh9Ty08wDCEw+euUJy0qoHZf
aGarxhePV+M7pPygV4F+ni1EtqSYbEssDZTlZeQ/ysm1ToyHwUnJ3v7uxyd6EzgwyN3JEHqNWNgo
Cd2NOAxo2FAw5oCWEWk5Xx6hIGyVh83MG1yj0gVfElNhO0hE8UYwW94TliXDUEe3uCItW+2IgpkN
Pq6WgIwKTiayZU+pW7kG3E9N5duvyVeXhD75ueGzLLFlB7Cod+j0xyhAM80ci5Gsyrmo7bKLB++n
wBhU+xgUrex2bXHT+xSPRJNhp5dXcn918hz3YUzoGHE6Gzi+eaS7VYAwp8YwVTWbT+yGBs2mxaOw
DwdhnRYJdWs1Q7HlTbfjWcMsU9G7ZDILKU/3uLAnLMk7xxU8YZ1yObQbCzmC4IYd6vP+ZqCcRrFE
1tGM80a5D0LKDHJoRC1eXp3JIAfvaPsFByjavAeIUe1UJ3Dog1W2IHlYHPeHZjdR7nHMabvk0wwX
OGowupSo+8hW32RzYMliQKfGK7BdAbpm+eaKQlr4txbe7Eg5qcmq89bRyYIxQvvprFMV51kR7pZ6
sMUlI/bjJnziHW/NS9r7v3yvdhSW3mvON4xNd6NEODZCAWWXUoR5ANKRBjSmstwJyLXKJO0Azr+D
y1HnE/hbq9CXFVU62rp35Wf8kGTD2M4g/UFw48J6L30y/oS3abH+b0YJDnmboPKNnXGid1fUYSnx
hHFabzQJGTquG8i1kIMhv4C6ngrkHVbZbUSHqFiYjxSA7w4p8Qwy7OQA5/uQCStv7+n5xcCCZiKk
6MqUrT4D64AEgggJjZLygEC0zCL1d2Fg3R+qbADxXetPjy+MAbi8Negz27ySbc0ojFOc0MARG/aR
Lobq7uJGaobJsJHHL+N7ypKvvUlausIzoB6CCtikFM1CJ+QABAYOCSgZu5k631zmSMhja227TaLx
8YgrPUHuEvpqcBlMdl7P4pkQFepspXNwBRswT4OgwZVbeD1WLuIlYq/8vMD0DEO4swK2gvbwhO7+
Kfafg+RbIVS/8n48OqFZvso88mYxPNFppIbW9OeUF6uZOzPDjMFwh0buxkjfyVP9n4olU3SGffv3
Y6Oq7Q26d1MKWBODQmyJ1+QjS5HNKxRRCniYbWHhwWnFF2yETHym5IqCpMiS6aXAbpr6iiqE0MMy
wnddcr3ROcaIW93pz63oqeM9VjpZQFXNBF0TXE4N65wrrFnb2+Z8srhnlxf8p1A1cN/2oE+KusUF
g0QiGc/4JcmqNuIYvMVey+SrFuppXKgQ6osmSX/zhmOQcWKki/QuSDYTWWQsAwTmXc54eOOauKjl
9Q6oNCkxrYn1TDf+t/1C1ncwSx/7b/9Hn+ARXcCyzZCHt3tnJK6Ui0k3LcFih8Lt+TBc9r/nJG+i
Ppk5tMxuUAv6zWhrZv7nYw632qoxgoICgoC3IFZUdXatO4PjDzWVXsYjUR+l3E65HPNW4Vcknq9y
l0YzwYX6vFTGgfCWCCqwnR4fjLGebcrdO8NvkgVwcU8IwzTjR7kbOGyttVPyUeQh0+0Jg5g/Gj7M
6oAM02/Qh9WvfIlEETJIRNDYkdgg3nz6WeJ70tafnOuhQs8Kvw02/6p2RmjpWRHJ+lezw1ABeUc9
uIt+NuzlaYA4DsayF/rYFd8F9jJ+jpu2xlumUGEhIhGjscwuHrPxEsYpn6KzEsK3hH8Y1T7lwuce
45RrO4P7bQ/pbSn4DJ06czf8vo5t2wJOtmLYwyAmfU5wAnv4ms0XNmtNw17niUAUfBRQoHcjDPw5
DNqc7YmWd+x9NDQ4X4+3wZzw0OZDmNQ2N+P0hm54OOPpLdcAVa6ORhnsGN+3vkyCbU9ACxK00yAh
blkZ1BAfa0jIny0wtlBqoovYKpvbdzvS+QsXO22fAPLkhV9THX25FtCkJ3sCpelNwQxWvKb2oBdX
GKOj1dRr029dGE1aLxNnhBbAKeDe0a5NxEHSDbRPsgadVyJW/5F5clm3XZ9PbknIKIZFdUHG6IXo
lBGLcZQpD5X1Hs9gg3e9Ww8uNmeAAxi9GGdhxDW6s2e8LFohXADRU/eB0JwXvwKSmYfRwvirnxuF
CuT9d1xGMOAM6fJmw5vZc1htuonZsCtDDvFtZUZqBc5titQQYNs/Zatn5OW20z+OlZkLuAfBdtzL
WWhlaIb5btDgPImqcqcoovY7AqpY7sz3Db02VDrNkvzgjkUuCVATCJDkbzK9hTtEnJRWY3ocYrHd
CXi7hFIRlQNJkpbNB8e5z1T8eNZcg0VrYDbvcFnLjjkpzpnes1bn5GaRLdt89PbSh3mLp91JZ0l+
gmpxpLne2f+3tWz6CgXrRLGr3uSisJwxK2CrFr8ikjfeFTl3Ew4v0S9ukQSNYN33K+QPnIQSg0f1
j9ykGNWfjERhCTMGavBQnU1ge+5HHuWPlHMVsvDgTYGbkbQT6NCH3I94GgG6Db9L9se+cp1I5XIq
9XFn6eAFqlDiQqMuU5LAFd/deMTeawOQbnS2HDETlOZ5H75AEvqc+hdfysAU03Dctf8jFMU2Wgoe
xvfUAQPHu1eeoFXvG7H+k0OYvAnCe19A+9om0crSXMi59Ed646cgYifsw1sWI0/pdPQI4Q/fxTRV
s/gJvytRhVnV1XP7v/S5ThJ+D9pQROvdej9AO9dWuHyTSyXxmF0j04BvskykAR6DsddVps88IMgb
ZdlrM1NBzaq0UAB13w+oX0XlcOpfUQub7ECzU3mbFVx733M9woKLmqbpEtKMVogZPXVqOJiA5etn
f2FWrdDVN/NA5k/nlxnNAe9uXnjSBSfytTbsssZaIFIpIVzFJHIBtnZu1Okq+0frRBbV8LTr1jM8
UGkApJKNI0eRKWlOhSqGI6MFKt0w2/qHValRDJvyFjxZQoXjr9jQOtLgONhVf41nxbvxzdJjErHC
+KNM/d9H3CaXw23kQJFFCN2qBcJnawfUKqIJHC2ySTqIwyaWlj6xutPT9PwOPMtXhvTnuFhbsRzS
TiP+DTlwaemOrTq92pvuVzohKsT169fVEu6fESb3oZm+r5pUjSzUNH+x9A4/yN++3BZXc4TsvyCf
jImLdiByOwtO7Yd6xx4iVSjRk2QgReU/TuJ7EjO7NXFDEw4oOWPy9fv9VX4ies8qyLGvj/B/i3YQ
BjKwrCDnn7PY/En6RBr36/L8Qa2OOk0b10dxHlvRNbFhrh1V2lqG+Mser2YJGX3G4MNAysNlm6G+
juEo1NLqVIaM5isuQymNzjExH/6ZYQoNqjgkNu7/mBZigNvjX4tdZ3fKs5XuASBxgOuleJRWxXqx
mt8l/JR2XORwURHzOpvHfDYIjy8Ib7YYrE8GXs0/0a+ldi71/OlrOxy0dwFd+VGva1x3SVPChRvp
8HONtF+nT7Rtum92dx3Rjmk3xaP6I0hyTZHzptPZKU7mq2QhRSSuiug8vuCGG/wM+rOXi9G+ZHoU
Ky6HJW6gZEVPwa+NGJYJ+QNXLoHXliAxqlrkagCizb5zeXQ9Q+6+jUPQimKWwLCb3C/GUEGOtqRO
ehKD6sQB1UNLCGhnD7c5nXwDZ2mITp6SBtwQMIO/rM+LAOqgVWQPyShivo7A9Hi5XLqUvpI/p5w/
Ux/W08oXpeV/70vOWKUmJiRVdotxP+uDr+cFbR5x6Bnw/J9ybcigXxdft5y/0UTKs8UD7MdsJx+h
EX6NlKl07xGHQrnfVJlk0TO4u1LaaVyfJW4P0kDcuIvkjfx0X+yrS9uhke7fIEUIioyCaCJxxVZv
0X9Bk6v+TicMG2r+q6e6Ccltshyp4UmmcNwrIMED8s5eD7WLMIczPyutBH6z1R7/Jscj4bhdd8nf
kEyFawt6n5RfDrE0WYuNh32pQy36/AixIolyszGIPg5sK1xXvQq7NirXk7xOceA+BrY0dJyq6aq9
kg64AJn5PYqY+X1ufpd8oA6lkhKjrp17ufsxwFKB6Dzc/5Z3pXFqPFAb+/IU5d3BQwOs7dfYvCAQ
j1beQSaY8fxkf6w+erbFbWRUA/smHWUqKCUjoK7+h3cuCnLe0SYrn2ByDcYJ5ddlDYdCBxWOPAvb
7NFJO975y2A1Gbz2p0YxuJtyCw0r8maoO6FSUcasPWdxqjzx2QHlh8bpRpfr1wDXwc/KDKYlfcxa
tjKxyJ2i3P+KDRcayi+q8yKryPM31wlDQnqc9m6SZON2RqTiXXRMggIfrBJpgy1vzTfugU2mu0lh
yKWcgUmCe8ydXqfhhUSOJf7M200v6lsPq3sE5gigUxaixjM8qn1DEIIEFmV6KHLXqRdl6tQ3+2SY
VNsmVIFRVTZnwWNZiYF0UrA/0vAINkJM0f4rkmgAKvNweatDSGGaSdXe6xypy0SjIGWdjQx4jE7D
AicqEsfNah6nkFDhGpOmypGDSjShT9HVwhD/Hu8yi11+VGtyRQW2cOZEX/bOqKbEt2S4u7eA9StD
6p7DqwEAv5er2m0XHucCks+gijOR4mWsjMMFZUVtB4F9Da1hXCaI5E80Y0mRq4mJ0QeXfbb8BL4a
b4d4sRzLc3KICmPmT06ZQvneSsEhjcVntuBzByc0ZAI4La7Ng09uECSBhHSqRSV2pEarGFPD2Vdg
1+CuArZ2qI3ewJV7j3/wvJS3J7rP0HmfhZwMCfK4okBaN374Mo7po+fGzbesiHV0ikwE1YkLn6h8
Bzkc17GR73dZVRJRvFJnvNLkv607o10uW0R5JyV7XwKIkl6jUVK6+Dcp5929xoQ/g/wV0Ai5EZAU
FdusUL2QnYxZCtCu1HN5FOFfWi4LIGmuzjdJwtkElwiLA8ULYBbmx/99eSwRwcmWJTQpwu3ysy63
3EHY8XUGsqOZy6o9Xbyt/ciCMnOknQ3P2gomstT4eSd/kvWQnqBOTHjvoV+3sMCmec5VI4DYbzU+
fjHEmM8Z7bRspwIatvXTcO0coC8CXSFngCKUKlXoX4VIOXHzzw5V92q1Ozq5+4qCM5ULaDg//jhx
W1qzOa1FVDID4+loiEV3fuKEjmDurlyilIDhvem8C8uqwz5z7SqWibgaYlHh9b+ZyHWb1pLqgy2I
LhiADB+NJ4u5TL6lKxSjwBVx7klovDiWUKqFbWqV55E4CIeTbLTsMzZcIVQMtgh2257tdGT+EEe8
aJCrnLX3sLvb1bRgXbptmpf/9b+KL0QBdtVbWzRzmbirNHaIXDP4N4e2XK5dz5ajNUo2NA07MpOs
0qGy6/8+Q1q8u9H3qaDbWh1nwH2Dfq+ZbNTWdstNeURKpnwp+e3EVbxCH0Mpmo/LoASznZ6m78h7
RqRepb6mxXXSOUV85AH0OQMom2LSuknvum3blYeiHtjT98uKn6k9iFPbAdoMombnStKB7JIsF26n
WJmYm6zV4LBnjFDU/Mie/a7MmK4okNPg0lsQ+7vSVNm9T5/M1z9tFa/li2otozy652ne6sKFnW1j
gHUWgWuJpfnd1u5AGIQGrVEnU11hg3IASd51S27Mp0UVZnrgiiOr6aD2EMBGwRfZaO/7fPQYYwJM
jmTuN4QbhN7LS01XJozTC9u7k/cQ6sNh1CnV+XE4gdRVbe9dnUShicwEEPQuKtJR0Jl3LD0BgvqW
6CpamlgJ/9ZFkfwrJOhmXqKNa1teGygpESEmP8eVY+WKSeFFfIOzDzog5Exx5R56dGkYTVQRxVu8
YnrphZpseuSdTEuZh9xYrrHG+vvNVfm06+6PiJUA6zlHbOo1sUWX8dLLkywFWp6vONNLFjeVuEI/
IAZRJOuyGiVevoSP6SOnDzeEdKWrWXFo5txk18sX5F/Lmfcz4uywWU3dwS9Zg/WEO7SBu7R7Bj5+
Tg8rDJrlTh9cq80xhcmfci9tmKl0suA087AbpPOPdHW0+F46a0BHUe5zl+xWH8oTj3ADEzvxRjBq
IDv8wb9ZGKvVSXskgB6vtaOAqtpIOks6V2wNvR308sDKao1haQ3PxQbG13e4gQyrHzyuhYi879Xg
1wdCK7vjQgALiFjElF8VTe0Yc/lTaLbI3dYpty3J2Zaw4O0V38pL5dicSDn6yUTPmm6/ay8s1RO4
Hm9Xyw0LPBio6G3NGFMsNMocDsdmRFE5swpRFYKgQBfG7wY5v5ytTP84rErlc2uiwlYy/Rc6RnuW
ovwv0M3JnlP6cJlCmo2SPTWb0VTNjtUgO1wk2Oj9cw7e++EXsJEEj2zokAdBmKZ0T68pJk3ka24a
+7L+BMGi9hzro2zWnOK4b8dKlUTDDcQIQ8ozJYyZFogJLOwfEKAg3bs9tkG0kiuGdw63QgPI5DWH
BbI/yhE74FxdPCuN6mFIbov5gUQ/7eabT8flJhf3yRCGxvnJur0ZrXnlFwwe7+j7H0rKCY7zNbIG
pxSTr7lv+E79EYEhMmOIlWTFocGElpncLC7EulClAXQCYEPRvjdIhpJEmmSB9DhiGw7J7mVAEItA
V+QZTr3EK2p6TGBF1zFcSjs2DtdprfbgQm74dvplUbZcLoOETvodvwIlXPe0p5zf7mnFhrTyVomg
BywEevES0+YNQpSS1CY2F5pYlLMYPuqtkoqdhUazN9r1SNBbVXXF7VJjFP7uTRGzsF8ukdEMHzTk
/dxSmGSl9kyiwjzh8EWAM9eRwYABPVh0ia1JeQ3nseP4yni53mpWm5fWX2QHA4ztWNZNJ8QwznJq
V+9+vj297lRfJvBrf62VidjYsYZxDQCTe4A8j9f5knjW+JBTgWCCwMIbm/9jT6w31CQ6VffR+XjF
UFOdt2VDUSIF/ssOtEeLlh7c/pHAbEaIcexBj6l33pViZg3MWUoaS28Gb5XhNoC+maN2DprE1vNm
younujv0CzV4E2fe5WQCVU9XeL3JJh7Qhmsk16oG5iGWjbZtrX/eC+xVivblPIf5W5a+dim5ECY4
Inuf6PmmrM/nE6irEJvG6oUvNLJX/yF7OR1K1j4Aegb9iBxz21jYK6/c3gKptTSxhGuvTEG1IjdK
x5ORLbBwfTuS7i+TgrwOrFL/zWtt5pTnqQGL7YdBdw5S/78zYqwtZorpv3h8pbPFi3sZhBxOTVoX
mWp+VyP+Lu+L4e5Lp72jeHe5JiF4N4XEdfR7LxYIrxguirs5QfPNljVIU1epjw8ynaJ5f82amyLx
c1ag4Ic0BuFdOV6Pqv3b6yMdCB7x7u4+5aqUE4+tJJBIu70CKA/vSM6nCGwJYGfeALN9e8bGa5yA
VgEcIEgNRe9LTiMCAs9sPjdoOzW0lpvkJ5TuL8H5w13TY5v0/kuz7zZnRAbRykxUGz0B88apj4uo
UHJtwGdeYvs3jdB6oBUp9bMffgFO9E6R/pyk27Ev2yWlMTYbn28nQFu3rs6jgp7PtHAtF7esL+iR
kTzuAgpW2C+q3gWqFgSrlLg38KTzg4gee1YFJxYp2F4c3cpzP9cE29ZzixM8yYIywYxiLHKEhA8R
OsIjsrrjvqNzX8W8a3EC3fDP4yCiShlxZjgJWA23wSqaxBXJ1qC57zy0gV8kdfnGDNxn9XFznBOB
lqOLiOqnm+dXvScV75B2iSdnPzjkpHzxF6C2a86ROD0i7vz+CcwLMK4cfP2Bk+yJtU2T8T3s1Vmx
Sw7RVVrm543wr0xxug0bccKIqatqFiEdwFx5wOQcoJVqwyASyHdihEzuIsGcRGvIhiNrNOMMY1sw
cn11OWv3EZS50Fvx3bc1Qv+5x1nPsl9TZy24iCWkWm0b5+v7HBWUhd1jnAN1QrpeiPY5cylNTX5P
BuNLDfEEmjbsQbUGB/fqB5I2/THT5K9RTbxFSIXx0LAI2weIcUyb23BzrHl1hYS+7yac0W3bXR+u
hi2jGx4Or0+HNn6wlI8rIBhWpUBPQmzkLTtAaX0dUjytcOgLH7nDOUP4JGSSD5M8M0ghctG3n1s2
kpMwImAL1Aqmj0bDuh0jYYyT3DhLxeNsjxUE4xkQPfa6YiwZUf9jlyV+xdXvEQOZdrBRG9TZtFpJ
8hDzjhCKUP60H+00DcpzV+U71WCaAtKT1SKozmyn5x+my19oLOv8/XJjk1OhJmlCcbOOdOKDL6jF
7sW15/QdMQ0K8iHcIJD2o5aFNBXmC1a6gl9G07AmvCrHBglBcYWArh/yAVCIlLM33XMjNCM3O9Nq
yE5IqLyJb4SgE9mR4KaJHb7sL56rEPNqAGy1l2zvWv+q3O7H0mFyeja1OufeuZKgCrtaHvm+DSwd
vb4dUDCnfJKvXaz1TO7XpPQG2ZlO1jfV1znUSOsL/DjNpZ6Yt8WtmdflHiywYTAW2UZcOtKumIg/
NjFP3a+00AyURnzSxuOWhLqXX5TUgPjfobaei+qCnK9tNgdPJIrAmowFmeYHIC8U7Npgd3Pbe5kv
6fOU/XNoCv2wy0qCZKI9gnm1oIXdR+ievgcGlN2JhpvhVIoHJipyTLe4SifvKjmpr7vv8aKRFXky
UWkpfi88SHI7vwlXvfO427XP0li2nW5aDfkaDEZw1zf1xuc5Qp0rDlewd9zda2mQLPieBuVPlwbZ
gmjaYj/P7elwOdMTwGBL9DJHTBTwUbcIe8CyzrNYzG4T2Cu8lnGY1+AGF/PepyuUplqYVKJkFmZG
LTqp7DPeYKJOSx7c6U9kj027VNMTNuFkpkB4r77AmaPMeaj8h1VPC1FRZuy+TsCXM7Huo4sSGoBq
OzPBXJyVpWu3wW5Q454OJjYr5BGRDpf1kg4M0Mg5qJvdXMnUQ1R6wZkykhNpLF12iZgZGOE02mN1
lw8wiVAcwG8D3WXOGi0HQYT9985awvZ/O4SI9U4/twQIlPjxRkHYzkxm/WSluNZSuKWg1vBlZT/V
e6Dsci1/POT6hMjtfZlPx2Y6jyK0nhZzXWKzrYIn8eFbYY0UtiGLNcfCtOa/prRmBAvSzkM8G6Rs
qzspNUvSzNd82l/TVR7r/CnX5iTqUa1dbFNeAVri4BFD7ekNfBxVwyMWnML+hgdqxs0yYiwgn/MM
Z0/MU1qr57MO3pwNjwzmo5q3OEw9eD5sSeOAcYPuJHJ7x065c+zPxpVzrFsuYICJRLk+l0GmyJQb
3yyOznth9ZEib2cvIAixZEYIBKXcd3dgzgnSOr8EdiOx5jGJmFKS9kRDhhRY75F/4/idSRDLvjxC
VEqMZdF1FoEe2ABEnsBfQ0S86y6co2kow5L/8ZZw+8lY45HD3a2D87mX0eUUV5U1WDIOj3bm7g9y
V6w3s4p6mru+qWC3RYghpUgjmqdwSgJLPNyh06vezb9WyTg/vzv2RfhxeRk/5IoipYzF2C5v81DR
UnnBI9DM6Y/EuTy7+V/uZzBey5FZdph/0qBxtkQJ4QZgRzduDNF+BM5yunO0QL2bdz1D8MvPy2qi
Bnx3VChxiLnAmvzidySFBcqJQkgEQFVI6VlEu32jUtXFAfRzNpY620t2VtuvF9iLT2EOwSeU7kIL
5u+FLrHYhgHtaMMR35CQdkfhowZM4boW47eUrz2vwUuaH0o/afIWglpZBjA67y9NvLbCPjtPi/lf
a9mEE78o7uliSOAxREIoygpN4LFtaTNljfd8672JOlaji7Cp6iEP7K6BXSWAoFX2S1/cBg3LL7JS
Bg4LLL6bejC9JRuf5Dir9Sv6Wn/OUygkuipQbhkbQq46pSg0N7CNKDIRuNJT7dzWyXXBaHcd7wKj
/UcwV3/dIrYl+6kH9w0H4Y+YSu3I2di+0xoxddUdw7SgerFNMwv8dd0JfatUReCvlQSApnpJtMAX
k5is7eADdOvLoHhU8jXGYYlcPGRBLUUzOkOAhMIjL0Bzhvd8QMYX5ghNN44bHtsNkHJcjAyd91sU
SaaYbLsT5BSZwu6n/gQEsZ9EeMY690visFml3NTYTuCMVzSXdIbjHaMY7WX2rlu1VEJzN/Jod+w+
BD0r842yO1nDhTxjaFqgUKjPIXm61aRHvSnHUxmn6Zjhiwx5RxEp8elBsZnEfalHE3RU49s2aXov
DxHlQkVxai2PX20+L+LEWc0stolIvl5E2QJ6ew6wjvSfXKBCjNyYlt9QnA4fgRjWYsoZVMRqXlgb
KDPNej0pWkSzpSjwqW8yNg3kaPBUXlbaymVJb/Ua59lXQuRThbJo0kkEatH19NGk9lxcpJd8djfJ
J6HVkqLX8VZ5KZ9b3EhNiKeuXJXGicsB/y3VWJRFbV3/wtP3CuZFyeRG9rVWR7dKzWRh0fiJuOlj
94eg3ki+H5M+tKqohMYcPxkq22iZQDpy7bUS5fRIWhek4+BlGRF4h6KGfrvILAjQTnATebbRrpmZ
sVaPxnbZsCHgDq7EP+x5s+FoF52vzbVlFCc6x4itu6sRBW+3fneIcGkW6ulcH4WWT3deZL7ZA3LZ
sYw5sqafgMGlKiu5q+myAVqW7EKtckgvxGM/tL/SZuhLUHPrYtBpotVevr6pGAxGEwRZX90Sk5TD
QkOH+G+PIykT/czYAY8bQTexOb8sGz/bc5qulbrbrbHG3bGXSwmDV7wQTlGzwCrJNGLJ0MufrGUZ
8DL9UbmI8MQvi6lID50DLUWVrdE7zAB3BQt/vStpacBjBmcabgtmB7UH4Fw7Sd4Rno9Ytc2TA4jn
WcB5YKygA4Q5OkedsbzJsXycgZkQ3p0LGHsSHrC6qW8JBg1KC9hbhwQVCbYq3YoGw1h4uH9cUuSu
jKYp+UquC7nK488nNHmB7DEa3hm1VA7ggIsRewDgXH+Soh1qyBk0NiQTgwhws/wMlxrc4WmRm9gs
11usbqq4LMLSpaOoMZNuZut/OnpPWXUbruGSe7Z8/M1y9xouYxT9hOmy/Q8zKc/GcV5v0aqzx6E6
tqYY2woE1ZE13KSPy6j1KvuNOrZQ2mksHUDCqGqMxuQcpiWRIRpoY7YJBS6e3PIP+PrsS42N1L+r
wIO+jASaGXYYmM7qN1MUp4Hdf/2KktmeTr7P7I3DmtMx4iT1FlG0E022p81VoKcrb5o1+kC6i53e
k+XaUahHcJkbliT4sVsu1Hv+k/Wl+Bb8fDNzdsM8FJSOSJX83WEqrtDLCWJnjlBOdmwTweLYQyrA
2xTiT2UoTHwvJszvE7OPHz64D1Tb+uPRAMuOCPE01gV7lOYaTGIlIEKZpAbfDdl940BFBb7fTBoO
yp+uDVRDtiBw3N/XdiGl5YS6aza+/Kd4GCN4jlWktKAIw1SrmhdJ+ehsHCBI7MdbnQwXXrhiq+f9
UURU7TNplyntv1p2KjeYTUYtncOOjs6SIuF9VAq29xAPv/8bJZuqsyvAj/FchZLWSKrBX062yvu+
xts9XKPXmZBgC7wclmC6qXPxSZoWZEnyGSMsCksNov1h22unsnLT2Pa2eBIPme5EscRdCzR/GUs5
fZy3ST22QOuP1oXkNaiOy/yJqkYE4GVzedhV0kTjYxPiGrV8qlaSxVcUV8evH6fvSwQrf60cwQvB
GKx/qal08ToWkmHnjLttEQtD+Yh8gpYuLEEMminUnjIgMc0VaBy2H3aSCp+SeJQoNQ4IdF+uZeXE
awTotohMyrRokLw32EpK1zPyhiBBeUIgxvsSTuOe8oDVk8NAGwR7Pr9IuAjGXubNk7pG8dDg3VND
dhPODe85Y7qpLCCMCWakEk6AgsecxOL6qUYn4UaXVH0GjopcQrggAmjt3GjjGFzzB9TpduvLlcXg
rARexXd9TExhw22jruwmnl/wjJldOMxeo5z2PDyikblNy+5EBgJJ8mCCLtMM4j3Al+tb1NGKYOYH
NbJxIYRbJUFIMs5PMh274OeAGk6ZHmJI0uGhMQawUYoC/o3EAygYvX8u6wCmcviALhXUI1PwkqDE
87zO8Qyhkb7sCZeldCGqwV0X1KTjaeMI5/QI0vABJr5XfRDX+DJ4ZOhUkmAZp1vv1TCH1Fqu45v2
rNrwSUIrkhuMNOi3UGuw+S2PYSKSP7i+VNtf6crfkyyHwEIH5Zr4Gwb2fA3If/21kRQ+M+x9p+I4
2gMCMkNWn7OJF9UOm+7tuMnKVzKdXpLnKmb8xCl8GU9CN97Yix94hQ4fC1RRDKfo4d7nIQW9yq/O
k6tqoTmiGVirON/Kdvcq5JKXt6Swm1H9aaQ0T/kIBIEpqQMKWvYqsWrTZwZBRNK0zDHgzLRQ0upq
0Fv+0MwG+cuejlHnBXg8pDCQut8a8kYss0GzJ/r3XjWpmDt4WX0lcOtfALB0zz7T7XX5iqgsw3Nf
3RJNbGyse+TW4sh51ReJGuXpDiM6u4i7pa/AxOEePcaVmr5CDufw1ru22sDvy+PAIPev0NWf/6Uw
dxXl1iE5pw40bg3DUNSuvyIflaNWsJkmCLwMrC38R65cU9e8+Z3JGmduny0iIxNFXKr6q9LxB+EN
EUrFqdYHG+y3nNbJOiM11SSZoKKDx2zpKjjXIrpqe9aoY2nwZg/z0XUid1vOB1uiYiycif9Vel64
b7uTF1Qkx4uAyHKcLHWStiROU0FVsMRpoAJyNfm7/aOw5RnFITDt8iLo+iVg+AbYE1/qjA4yJ7/A
VemDW9oujs8jEahPBq8o1OAoYQo69nGdIQwpbEU6RQru5jagadYUgG/S/0wOOvRTFggpLP6oHGju
IU9369yfJLVTzBfbTOpkRRxRUBQfEWALmGjiN+zLlf/nOfn1NFkONOWLD1APiCUd04FUY9+6k+9b
4ioYYidfZZpR/YnKkaP5ivrAHF5SF+Cu01pbWCKamQMmkXSJ+qxj+/zEJz+5K1UJp5NpPIAQ+flb
Y6c0AiIzQThXsF7Sbimkjc69z33BZ53ZSZeP9SmKhIa12GoSgaAN9b/OwFS+OHCEm21UAAQRIEN+
v27x12xjkUKrburbY6rJK+pQNtxXuKcOwB2XvzSgn6wgNEjI+ZITFJ+c/Xwy3s6UIcE8YePxtnUE
pVGIGNUDVj8tYJU/7nColIIbJkUvwHrM1kOIlcFxE8mzpprl43nooBfL6Ag2iL/ugMGXgR/vzwky
Bdwp0dKsS/d8rxhli2xgoLufcec9KL86SMHyEqG6yLT/if2nJnKrw1UNMrqKnM9azAHCPdqIcfIg
9KohTSZMJ+FTwrvztINJavX49Dn0lPad0mbrZQO67XztXyqoXUzTLJGWWTLsPjwOIa2zGV8/pZil
WNCLkcxOxODVYH3GvaIIctW7n+EyzOzX0m7BB/hMqUUbYfolTqUukcra2TexWIA/b6BFDQZT6tNw
z9VwEtEUwolK63GfyQbbkg3NjNhftMYZmKuudXR3HRjpQScVMfJveDl11bxdbrZ2esszo3yK+tXr
wSH2PErjN4C1PlqwYv7wDVPDx4X1ZyMhbN7XcJeQbPe0/6KVosr8eAIv/z+BbXHG92QFlleB3C2p
gACMJAic/19xWTCoBdRUYElKMzutS5EfmGefXSHLdh9ZjoXlusDVAnd+sj2tKWlqbYL4LseSkSo2
TX+cXjm6sMw/YFXJbp2O6X3CO3DEY6REo5dUaEiPfNkar298yOMLecrob7Ce3QL4CtYOHmyWBS8S
4GPIh6G52l+SksO7l7yW9F3qO4FCEZO9qhuW1XEXO/qlGnFH7iQy7fCBUKu2nmmjcDxw136ysA2s
ylxFWyTzftYb4uNxc1ltwno+WLr20uKNCOxChCQdAcSQtOm9oJVPihaRXg/kcyBNjF2TmnJpVHKo
LWtOgkJttrWuHOEC/+rN7fnlnlQd6+UYQFCT/SkL3y60HThVnBHFMiqqH1HtyuxAW3Bhl2iuBC2p
QltTs2slZh4CDDZE8AYEkEgjXSCt+9TKtiLo/qXjEiVW4XOrdwiCTaUVn/+bOo0rrrFDZcMHbDwF
6NihlyXmkuSuKwgmM8Axa6DfLDhyIzvJZInbbLXQ37p4SMeA0tNzMAykKZcUivN+3NsGgDUbTPr2
n3hssDovxWV4btEOB8ycMxnB3Tvp9KyEZU5ZpxN9c1BeihT3k4V3pmGticCsMkViC0IIS6h8DRZ5
pyGsXxX8abWswDSN6SY0aM0tLuvjS5+fBoE+39l/tYxOPCEjla846Db5UJJHSikyHGEqvEBcmkHv
se8qnyMYwYgze0JmdXTx3Kf/FGPqv3b3jjrZslG/oKxOSqZPLhM2XENP4YBMr69ZbG8AMEjRFySK
VjLK/6y9jtvikNQ2j9FpOjPScQAfuznAG8/Fg0OG/4R1rM0eA2boTsKLTrWA89p5/2M1idUkdsGj
RCxSPTTGB6JwswLj+SXJfGk/I4OwYm93puenMQ7D/f6yC4O+eBScNcyrtQ7jWbtmQz5KY+P2EMcB
608w9TEZMXJ9V0RTdpAF7ZSeXIkC9EvxNed73TopXgMUF/ABVgaI18F6EEzUaABZx5vHLG76obun
7+fes+T9ic+P9tTzx4HT4DfrDcMRlcani2eYhW4YlqClLaEMiana2h8QAaepRWtFj4xE3loqWw7K
RhDMRY6NUc82eeCZNCU+0Gurcfyp3oNmD/RAnY1JVuvyw8sXAY3ydHiDrEcxLVo4hF8sUQ7XGtGJ
8j70uyv/U/21oieqDmQmU/xpROc4zjAKlEhdGjPt/TqbBu0ItohiqaDPEghS2j2dARiWl2Q7jAok
oRfiDvDTgtSbxzueBp1yf84wAAcs/YB8sQid710QRhmTGnGappomTD2UiFhsBu2QmX563+9zWv6E
P39oOwOvjT3V3tH1sHAAKvIwvnLzMQe8YhPqw14KtKaza0ymM7frQmdyBiYiNA8QHTEdQG877d+1
j2lsxdKotxVufpiEkbWTfJzQ6Nk/LfLGBOouSLvOqBlyYmgh66xb0Z4bwE4LiasHVXWu9W+ShOfa
4Jt1A2bT5J7QtDmBPaIv+jyyBu05fkr20tfnHUDpqyXNga07B6LE7lkymv+vvB+LFrJU3s4dMVMk
5eYmtjNpEP3tQLwJOVdM+v+3JUNFTA+xeGuQ1mihXP/yoL8mEwv8YGeSC43UHfaEZM2vUoHCbpNm
BShq1o2WJhLAfjxOXqo5LYk8920yGQ6hA2AFE1f62mW7iAl9uinTjavFS34LqNa1dTyiJwaxzxFU
3e6ASeI8qITKK9vtU8V5W52Es1EaqXJSlzl9yVoVdKp7g+xM7myVQJKCf2evPGHGCzeLiUBdHED4
/O/SWFBUQMaBRiXtiJ6OHnmCn8twdyllMn/GY73aSH7NfvRwF+sxe7nbS0gnSNUAF3IclfNkDNwI
5LSZUSFTrXS0C7kGsSwq5veKJokK2CDtCXEcTIR9qdLs1RKKgBx+NLPhO/SAljNNQLpRYlfsKRft
RHTTfz6cG0BCPzPTgErpnvwPeetMzs0/G9LH33cZyvXRzw2JKuZb9+4PrZEjwbRAMl/0V0bHsYFW
eoe7JIc4Y19L8+pwoTnVC18skBE8TzidKl9MoWKz0YNCPmbT+r5dMWVP2vz0UhccHRHn/bnxBnzh
end1XkFSTwUJejXdB649nh9pC23gSx27rHrdZap9FL7A5UXOAMZtA21KrZxtHkmtUYPZbst7+maG
ER0X1UdKinyx8pX+ucP0zWaCk2RbXsAk3FJpfjwDzEgij6qrfIDzJ19i6JzaiYndIz+wqT1yX3b+
RHjw1qaVdomLMovX8TkdAtA5Ud8+ig1qC2/A1sTiFTvOBC4Qhdi2KhZ55YrXGxSul/rvI17g7zxw
QkJcerVUggcHc+ZyMJjeSKixj9O7mhM1Zagv6mPDOU78OqqMfLVxWF5uDmn0qjXLspubrwtIGurp
npUlvNBZqvW49H/2NA2XktJW54XRgqAOrDOlCi/8FsXnxGNspW9/9L7gk8NUd8pw1bbGetrnHI3r
OXMTaM2BEb7gvy7UJ+LPwY/Tf+TCtE4qb9a4VRAcVuBORVJapwM6zkdhwPlWaHy9eFnkzxCguCuE
MMKXvGSUAXmL1lhs9kUnLstm/2qfOFNecrRwnfCGEWM77YUXuDLoQZ6JlwC21C0dJPQlR9LCUCJe
XHvgXo4rwwhW6G3Lpdex8hGlTiJzTNkDvLevFVyMx6Febw8UILHTCBkwQp72WjLwniN1qm+J6dGo
9ozB8I6FkqYUY/FiY5QgN3AMQROmdbrzX6Rqo6tiEPKJI/cCcr0PRWMG1fIQj7gAFeixb7AmUBos
uEhZ+DM3dk9g8F2DojKKUKGqVRCAAw/U6DmzFDsu7vsW+iBbVaBfOYGNBdLKqCrt1L5/KSQYe3cr
NOByJ7wYCXfH9IPYp5Rs9WKCxXn5Ncx12G7Nu52vfmV6j+yjg8QN/UiJEXnapH+UgsJjQL8K+K0F
GzfzHpRs651IjqbIStBehlz9z7ZkUb1DNUr8tDqfpnHSo2zIJuQyqvklNfwQL6hyntVjLZ6PxW34
eTatiPKmuxrfUrXY3jcPhQ6STu268Bs/h6i7cPG1d3KqLuxTAdg/+gTxSpKI91jXPprINFALK+GJ
t4ktnsvqadmqr59iUb1o5bG5G/B7FCZhT0g7PZRAWrZXtip4QMVFp4AoBH6m0cBWkVV5GPSs5pOj
95kv89RxekPuJq8gu0cfE9a++oQ1BIBs4dU9htdM6WGl9zZmU1jikSpmqlJ+IVdaV2GnO4u1kCfv
R1OUE7UzwrnGYsjNLve2GcOX9YGDNM6YFONabPL/ID5KddzOZBa88Fd1iL2xyUFwdcCwyeR84thJ
vZOR3551dQj4hd5ao8oogYdmeiLoGu2SnWm8QNTOGIlr2aWvlkvYP/b+jEbib7lbTCpmDcZgYxYg
zxNb1ScBPcONQjx+RGMyQQsVoxaiaJnjyfm10+NqZgt3J5ah5/+uzEiGe0LjAiwP3exAVL1jN9Hf
pFkCoTdUQMJ1BKY5lCNaqnBNnVoc0J9N0xeBFqmsKL0befpYYslFNrvOjaZPsaeyBbPixxrJ8YYv
r4hAeP/3yTtHn5iaGwbcHbDVZGeF3YPTV6uNntZy2CYaKJwPqaQGdDQzbxslzSNzXcfEIqURLH1V
FCqR4oGmhIKLE6wdjHIxsg003Dkbl0P4XLaSRVqPppFrMS5NpRCPEfiwoULIyY/2RVhM4a5/VyeM
kNusbVFAvX2yJb127k4alDqUB78n2PRPJcB7s4ub+hRK8h/BHNgIbIxKY1poIlOtv9qLwnvrC9e+
pK4BYYNS9qXwOndsftgNKlEZyQeOTx+SvhNAen/XgMb5wMlH9RF3fE754c+Uev/4ieGoPhlSBnBV
w2GGiBjgQ94oa+JmZnilOnMeI0DXK0bpeMhoTOLcvFGurKms+AENVKved//9uJyihx9WBHm7fgiA
+y4jrJLEpLHd3a/xwB80SnGVduUUClrz/XOnXUMOhyPHll0b50cGGi8GedRbaTDf2v5lHlZUp+pa
H/itbu5m9FQMQh5vPacj9N5lHBx25nWkkuMwR0/Z+O8GPrzAn2YamYbCMHBj2R2RP/0LaffGfxKy
o631hD6S4jGHb6niaE7hWtknILNQ4hG19mayPsrY1j9ecODryS56UwwpMR7mY/lSYBpIuhlrNgfn
DGa2wE+OK/9wF8XB+yKtDzCbjBPcgzDZ0MKVbYgzKmBh41maeNOH226xL6mxOeJpFg9HE13duQLL
BoEEhxXMXMTo6mdY8Ql+YLOO7MLju/P07l4xrNeLD/AUyqxQtNzJBLtoNZpuBq/SF50iVCcmsLzk
hUxdAjsOWjNfO+7ngTJAgRYkU0aCfHUAMBN/kgHNLrBdShtLD/s0rRvaZyGZxk/zRjw8yoKC6gcY
CsTZu2eqtXZ79SY5KqboS4M9JA+Q8lKGSCkeQ53Irvv38eBKGukzvyMJo60BI6CyUIVqcztvmrIK
dgogPQF7QTMDBpIn1yZXHaWAKLFwLHTMAbgZmX/Ro31asKaZShxdsRTs+qXNqAlc4qJLRZXBJLqN
3KBG5YCy8zcR+EO3SmLkKWW/RJN66xXToueANkATLVMW7F7TRQv4sk3BBDf3Y6yDc2JaijFantFG
xDhEqqlKdXVb6IBg6K71Tf71L8V87JOrb+to1y6gPgPXEl4E+VDfd3QqZvmfKefPhDk9onXMu7DQ
DBphLvE9meRtpMKVI8YJZvewTAWvnvTRZsECEHYDY3jqns5HR9lpzeT9lCzvyMehkp+OHAHU6Aa9
mWJSHoVTuFlItB/GM6CAY0Uu7hY4eslSTR5StEKVvjLyyA5idck+gZKy2TWxnXIi2gOPau9jvc3d
En/5dYDQWPz+P/xBk7ZWXzL0wqgqHoosoDALYAmMWItFzujfq7t80gB5XJFpY8IbfvIASUhE3kg2
FZFxc0R6Nnt/Mf31VR8N7ajjWQgC3s/s7BqLeEoafLIffhqsDDMdI2b+pc+TfI99QtFue1GGW9yv
Dydbff35U96laeenmlcnT0d1yRFZf/91V0qz1ogOcVNTUYwNOtaTAKJNJFJFng6gvBmA2LujWqN8
2TQ44Uu7Fr3+NWAzGoMfrHT77N95yrPEEOCd9SEbCW8Co+tKhE84FBBrqx1vkT+7Z7hDumyXLhvk
CY03pMKLWoYnhadnbOJ/01C75nE3qfcigELYTICjNFVD1keqUCyFNjJaJlUZmhKtbnNPoQ4KmJBc
yQqzUVMZG7sRbyxxxp4Zzkm0mrrydecDrpz6zQOuHHQeqyFTOxCTiLsTKsAroZgBdixg4XHoiv7/
hULiDTk8Nmh6sD2w23RUJJPNxfXOBU4AbNSpFiHVW/EQEWfRkGtSNOqQ/diskmN9Xmbke/+FDrDm
552wsa6DcfQwzwlPzXKmRvoOEyxoNPeNCjRMmb6SM1A5u+GnQhDHxsZcmXneRekQ3T+8XtJdZLri
+yqxFJqHnnBVbsM51ctVDkENfTBDh+AnDEIqPvjt2kdXl92PWqlS+yAsgUQDJyiQ7K8+x+dTF6m1
SwWz6SJaCHShYhbpZtrPrDjkqVxZIuTQBFJA0OKUHI4f4I2A1bp79tg5UgXbrjfeo4jJQlhj7uYb
F+oQv6RaOBAN8VUFuIYBe7QbXlGnZqkYWcBybz/wuIQ699XTEf5LNjIHUib7cfwuShdWh7EBsuVB
x/VZixNDVkLct/DuX5kMXlcoEEIz1yGxZslb6WVuphxVOPxozMoAYuw2vdVxJw+ux2CKXjIicYUi
GmBiivXKzg9mWWcdUE92GGBhwFhE850+dlnYH77mcmjekoI62+b8aMJugYdHP88NraizYlcas9Du
3znFTL1Z+8enHKO31zyGEC6knvJ3u+q3fewCP/JAz6Sfy6cMwyJrtmlTWDw5ieFLw4+SA5md37ai
PzpN9nfFcj2RjxANHotWhx08QWFBc61s+vUTgH9+VgjMtr8HUn5itkcCSuzScM2YTEwZEdI75iLc
+yTyNFEwWPdwqugzOphXWiUgy4ZMSKKFvy0QdPiaPI6VKF44jInm42BzbVArMDBIcO9Q8EGOjFLD
EU/khHpiMSg7BoXmBZNDXRASUJjmptTpSw0C8iHfrxOjksSDzaJ3UpxFkV4N6zsoucM0c8e3Ho9P
qpMwyb6PxK/nGhJYmvqYnzq56A9TyO1jofQyi6cCXY/17hMOoSXbNgye8bUSLR/gAeUvFEUawB3B
mDaLrtQMsp4vHJTUfFrlc233ZOQxem6MrkN4TUYP5pgrERuWrR0+pzt1nFsVJBdPj2qDMj9OUgwN
JA4R8z951s8tjbQA9zlnZ6ei7EKoAcavJdeqepe9yTWTPlJeKUhF1forqJs7HkmGtOBvWJ8eFm4B
wuTE+q0McHbMsCivHaE0ZEua/o9CX7fP51qq/j+vMSUyhL8hV2BBM6/H7AAUhrs0MQ18mdp6sZJN
106bo00gkGau/4ZpqQHIudEILPQZeerMWJBvY22sPrATo7XxBLJ4mwxoD6uvEOyOdaU9qH1UpZOQ
TUK2BBKEQjaw3E/d+a6J42KWrTH4Ac/Oxe3xKbA9DEM+7NFciv+5JjcutiLwfpu6r7jJKwBWzhVy
ZpvP9EkLtUJiK97A/EraAovyk/SEp2hXloKbqOJjd9y5mwYVSgVpS/f6ZB/jDkxpWnprozg2fMA2
STaOYpmVvp2mWiOLAiD3AfIwcIuPUBeQcm05/KQu0qzi0zHLwyIaJdQAXf9o+dNdl+S2Ph9P4Els
Lvge0JshUTezitHryRa/ZAw9E8NnLv3AtVMN2WCHPdOxV2Tme7cY1rv3sjSiD85dSHfTbUJWBNYh
FRsDjPkqXTWVPYXEhNikAVuQUCPl5MIEGUjuHSWczNulPMQjZcH6oOqER/rEnBhwJHv/Fxp1Wl+z
7pKLdUip+ZGdB5GAt+79pSkUisDo62ZduTSgUi9E/0SfdjRgabWwE2zfghp6V4EqYgLbBLeWEkLy
hLMb9J9NLhJsbOz6J36r0mUkqZsa1hokL6f9rCne2xHYOd+v7k8vzjSSioH9Ii4yu0ZTL1FtnaUg
XowqF3ZIx4cSv1dviAVGBqlp3pVa4QWXXGpw7i7OzjgQi8b76ZH8JOH9BRwKcDf1thzR0ZWKHWur
bPP3JQyxsgqyqM+8dJqUwiOB7qWPHaf/PqaUXTyDQiYEw9svUanqXMdNT7famh87eu+3Lu2Y0+mA
3CH6A/U49NIxjWEvF81fHmMjHcIgg48XBwycNvV/6Ij5eDZc42nXIUwVRwALiHu61XIIvCFkN75w
N/g4xYkAmvMsmAx7wZtehbfHWTH5gFNO1FFyq6jttpOTOzEDhuC1dpCkw3SSds9Smwkru29jgdO9
fg3nK4S6h0yG5GKAMK+AubaavzIzLPX+1u639wjR4O0KZSlVoKjI3x0tdShx9KpbXMcbIA3vEkoJ
oSrWjkU55qNYHjeVInfo9zS6GKjgAprfQ5EAPE3yw/IeMVR0/fKHRGyZ9ARv4m83Xcqjf+m9J9d7
MCCGfIMLlTyOJP+f3GU4eipLWeiWW6xQo0hfcuCBr1dSvZKF5TkUh1dfJsFCsTwbD7ydtQ86dwci
7bkFV5iSqdUevPpBBI20IODlX0lNFae+Eb46SDd1INgkt/ur/pZHApS/Q48nwKUjL7ydhqs+KZRQ
2lhb/N8VcBax2xWYrZVYZy5YV+wQ+6uRv77y/EjynSTPcLDVBWuiljCEGh1JAyoe4sNtO4Mq78cj
JIIvlgH27HbGzjAzg3n/L825ZvmWBAl9FI1rtn1KdgZIIH2G214eCcRJQU0LmkrzXIPkwRBUL4aM
M61XHaR6NYpjfSdv8Q+hzf5J2EmmyvY6m2EqHrDkwO7hl2apltcWzXpAAqckM7YxXz68PzJyOSDf
ZhJ2KhBh2NoHs0uhqnnBXiSo4GAOpm0Ua2PCVK/UERXuFJ6vq0FXxG5jZprQmlQhLbcwndfrdz5A
GofRpOY4vSa9Ht/RgDMS43Mqz6fQ6BbQZesDjzEYUaLd60CimmtLCVXxWky2FjfRYd/SS9BotDV6
SugHROMZe056DBabuqt8p9en0e5JOqp55yZ9/QR6YM3m81aNOFyTUlJ26wohloCrsSQOYUjOubeZ
a66QRK7x8KXf2RS0w+gwZW5orw0Pf0ss9EW1OtS7mcJdFIvEEZrTrvm9jWHcoJIsHqqS7/gqxHla
NVu6rtLMQxcCU9l9unw73JCDaG7Ee54j39mFAqzBrPj4NlgtEGbmj7T/nrMPNzyk1Nr9A5IzSP/A
s3VXH8matGxRcjKjrlQw8CDSXZPsqVLX/xrqJAq003W3a52qU0F8WAYBAhx4GELdSeMbjpLPqyI3
Obo3EYiMzTYFo5fqXvnHnl0FTuuvXRU2jKWxWFX2M7t6bj2AKtdxrx75bxTBETcv6CJkOhuJ2onJ
Rr1oZhtIdZdPGfnb50PSvKgD6a3/0u5nK0b/kfmJiqAi7Rdro7hKOXVBTCtWepVUuCK4EdQ5KphX
4VjdTOxANU4NE4PM0oEBlQEzuc7gn9qTjYmITK7MUyOouMO+VKzAsHg5otP30iNvuJXod69ZdvZ7
CtGXN3SRnsn1dZxvnaOd4VzyHoOC8qpZvKkFpwYcVEfg5i/SCARWl5exDqaPbYULhObD0axz3ty4
cRbHsMdvO1wctvkIa6/r3/gqsmw7PaLgW8Ipyc4LdMx5YQlovZs0HXBCavQnAEc0/3VCSeEoAdG/
gkYn20sFDoxG2/p4eFxGhVUzo8LsQlb0SKFymEaMZ5dI/ZWVce5iIY8e78geTMi4VOj5RPhMoTDx
WfGZImDNTfb01YshPbJefSe+gJh/pP/mlsz/qI0kVhGQQ4EANJw9uPwDx2t9dRB8yWNM7IHAR36g
9Bqp+Bjx0rdbr+rt+cPkfVEcNLnbA/Dkpn1TDj03dtMkMJV8kU4dyBjuM/lxDVuGf3/CEdBv3MMZ
t5o/OHMvWClSkT2SKMnefx6EmaLdzpR2h/6GkgtBrRTrcy/fgVKI8Pc5COPQVEZuOXfGyWdc5kS2
QyUm3W3db4f9jXjfROR9037nSc9uIG8K8rgB4MYSXYqPVRR2cX6hy0E97oj6wV05CMyfZJhUsuMb
5NfvLABr/N21PQOCWakU27A/1Ibbs7AuNI0iiOQ3v+D7IcizEJY9iK/ekrEBz1VJjaoDHC1FCLpN
ZgaPdprrvtuXFEzwFi8Ph0TA8AfGAv540lg4lVYBlEul7b45kay3mNp2pVIe3OK1CzDOhqkrY3uI
zFZaZCIPiCq5sgJXb4LndXdEl0cEmh2akwc2W2u5hJfMtWrU0iKkaDXuP+zavZ5/S+VSsv2els66
LkmL6G3yle1ApupyqEhIXJbAb8vpkT4zDy4o76nLHusqT1vUx87XLPuY9ANPee8GcqbPOaQ/SSma
fsUENpuchRi2LwL2xF7XoxAmut0n2AuktBoakYfG17ZZqu2LEGw0bewsTDx/je+KQ82cgVC6Z/Mz
YaG8v2y412nOYaVl/zXSxU+vSoS+1cJqrdm9ALyoPvpdyrnMh6e9wYbArffu7NbltboCJh0Cd/0r
ViwtpHift4j7hri8cE28IjOGH07eErKDYd8Y+Por8bU1uxhhLu9GarSGPyv+IJpfsJH6ApoEyN8S
NnSYoYyLhbFZ9rmQAHBTDQQeaImFWcUayqlIpjozLXW0Q86NwIHoIzGFGj1gnjq/1eub9BB73pME
EoO4dQIIQSStsDwu2w9IKaIIUVWjFB8e+98eG2bH7z1JjmBwRX6/lof9UTVs2olk0O+WYtPVucfP
oO8oPxeV5Eq4dE3G9fTCcOugGMSKOLAYJm/3hcygQSBKOytqIZYtzakVuXVN//pVZpIcC3h6XxZh
303ESBwTdpU7BaWC90ALYrSf/KnAS68GZ0xA+a0II53VaDsoIXE9NEOhuhPJ4Rq8G7ivOes5pg7x
9eABz8kITo5l3cpc+gmCGg3CFuk++NwrOqW6sM6HDu9tGKAqVTZQmYvpPfUJVaV8IKJlCwJwA29G
SS6YDq2QoaPgQ3CwVZSbwC/qsSRwqqxyLC16HsYHlnHrFgreph2Hm/bgb/M7uXZz1f0mEBUs4xsl
n7gUVl+O9aORG0E+Wym+0D7KMWNZq5QOKIW+QZVw3EBChWpK2mxhxZkGLFSbgywoYy4D0IfFjXCu
r8xkdxutQw8jHkmNoR4Lf7IwXfpjHr/eOM1OzCiGsJPWq2luPID6Gxn1gmn3rRtZq3GPJ9phWVIo
ae09gXmhHqvcG1USQDaMhl3RVIV2+3+vOhrfBeIxBF1rE27f4YIRplJ8u2wSx26bhZlF0i58fJ6m
8kAOV7+ps4owhksJEQG3G8aSfyJMFTD0BPHE1tVI2JWZq8YqXhWJndHX/W/gbtHzcLmCMKLCaDB6
P4PPGd+U7JTcCaT8/r0BrQRSC0Paf01vI+Jl/u1STjPoNHb68bTMtBlAXRCq6zVVKHDho4DSulZA
D5UVSjodkQWuSzphI0Hi3mlMmfwoKhz0Ny8nF8I8bM/NGS9SD3Iy3fv8QkoBAya7/AQL6G51+lPa
ITCnR3v123uhiKZpIjKJfSUd/5jeXdmsa8yA98nJBiQU+IHvr0y6os0RGcEFVjGw2tJBA4k+xJSc
PqDor3IS58oPzlQJn2YLDgpZyUTcWSbb2UzJ7YhbhZg30513bEhI1mPs9sku/J4Kdq0rk2dTgJsx
X9trDpnYMKCJXTADDu66o8gTysDEACS9dOIt7Xl7V7dazuYF7en6v4WHUUYAdbiuzssVktbPRQpu
mLFxZ/MkWNCJrhXqzrl7FZ8P4hEQ/ErrFuXzd3wr/koszMre0WV75R8mjFPI75Fq14SGAM+BzyFw
HHQGFks8w7acJskOzrDUwxf1zR/XbLbVSMC7RdqHMflU478GDR9RQnBoV3IwRcJPXECLRnXM9r8g
J7PzMvrxj+bVsmpCNKy2V1WDszcH0vmarlsUEPA9s9Z8piiwTjk16dTRjALMmwCfbiM3ASU5/j7K
2UJRu8WI2FPyEBReDEriGfA6VmBzKEj60rcwXiiup3jWxGj5SrsRApwiRaSBXOATfeH4asuofTzA
tC0e7WMTUj0iMdJ9jnPHhzh0qtDtTKv5izsPYV7JwuXWL4kLtti69qwlFN4sIaSax6nHU+frB2le
1rl9dSXSZXtoAh+mGyfd+QsMNdnkkAzRMEf3xNDJYKOVFc6VtRebT7RHv7gZkkFu6rC4Fu0upNjV
QxB8QpSB2jPk/CC1sO2stl2iPzFKQ4B0ygoKB4ZmD84P8EFQFYTwoi8kajkucQsKYLTxJDHhKoow
ttJLQMiQRWdH1pK9BAbEob3+eJV6ZTM2UvdrrtB6wsaNSZ4JAalJfe4GxKDzq239cNKqptOKqbgw
kDYStWT09ItelyAMQjZzL0OaUnAkA1tepOvv0jYcs+Vdg47RBcU8OeFW0EbVtkcKZW/oni6YfFcV
JgVsBZyUDRR1soQM00srIHOmkEzXGcnxS22veEfqA5KiZQkM/bAqWCYS1/kBuc0zp63/FfuAv31S
o4rN2/cuzzpe/kpjJ7qg3ilzuF0dVqfMQKPYi8UlOynBV1y+ASyUoXyuZyHV6wy2JxGWIZkg4RUB
dDXkRQ2sPJ2S40CoMI/KcCHODsJzNu8pCyG2hKiiHuOaPIjQzVGIZOVYqnsDmtWlvw4Nhcs3LxdY
OOaHDLddU7TAnz1+no9DjvXsDMwt+HMGRrWH9z1WejXl5t2aqnnC+t4NoJ7fpylQCSR5aSq+G/KA
B/MRUsiXmDhyV8qZsjlelSBKO9x2Lu0wad0KSkKmLbG9/BMHj5D4l/exaq8J+8FD+EfkhbK+p1EM
MVb5zlTHP+DYKyUqbSjiwv0k0AMGqA1n+l3mnoM0+fzgtYLXaZo9V/zzXwpVmTkLvrZ4+Vknorax
EqE6K6olSNBNjqYeN4UuiKeh/q2mPMJROjuD++A/njICvG738WMz1EAvxzQy4X1jVjcXZWpcHiP2
wEAaQCbK4cVCWSWZI1bGZ90SUCC+wTfy9S0ahzyEljU1xsIGTDtA10IVgNvS69WMBc4KIXTuS2P3
DE3ifwmVD0vj1XaZA/GQEcgVdwKoiZlUodRIzM479LebFQYxChRBywIlIyj+kAfdwFS5Bdxva0BS
0ONxRb0kdEhLXoa/6B480uB37IVXXhECvKi766ZOltVs0HgdNM38vaq5aexkZbIE/G140Dyp57IU
S3ybXbAZ3Z+FA8zrfhrTJM6xmfpchQ4OO3BgVEEogMr+ksVSx/katQpFrMFncdo8q/kPy1bPopbt
m7HD/sBRIadpPFWvub2rwHYJQkh944M7/qBBw3yKHDrmJPm8bw8JyzkYlSZXoq3r2GskWt8jxNbh
JT5RJYJljgJ4OQMx1ECei+wlNPgw6vIqsz/qdg6DyGxSTt51IwjGGwVVq596Pg2rCBmJg5wSxHqk
RZDEWyWfGT0pmm73H0bMdnksU3pgKiaVkk1kyEfex3k6NBJDid2RHeTcvlEyeBE68xp/AT4EnMTy
S7+2PE07dJtjkXeJuq3MGHvem2yJwStQKiCMGFyIkAvgXIYdlPCgszg8Duix/vL85cWQN9E/zm39
Pej74pLQZGoyokne1mfCuwqhWkPOq6R6Qt8uYFycg5KHeD4KPqyGkmZcUyoD2NHCqc0PVTSF+6HW
bJjsB51zxYEasJQj45bF1lp9BOwcX/Y50FbxxC7nZC4wVPoZlBgtuYKGxkM+/HNBF32AAs12fJQ0
xXjOiAbsj8v3WbA4ANZh/zjI8tmNXYFdgpIJ/cDOkxkj1kYyYzxZi3qd6K2wLqLWkKbJXBrUqhv4
1tghncyb6BxbA71lwK5qhsZHDK4b1W5cMdDZfYkkIxqkS9tFDm0enH1EatnKzjAB03oS1iDD800s
X8zxyrXm556ydbr4bHyNZyt2OD7SNithWF4NtRw5tzQykTp7QpFfqTiXOR2OMG2QfxZE4n+aGHQx
O016pZ/2wJkB5EL16bokEN2qeV92CIDqZahIJvBKO2Z6qGEUiVjKXQxaWDmVDA1WyBlUFUspchz4
oexGOXAUy3ypA8+j8rQefAXmafAt5OXZlIy7gQLGF0bn+/YCCfWnSN5fmLN0VCf8WecnGsWGXoZs
7Buy9l5opQDPqgkMSjHlqQmrpLLUHgScnM3gJ2bxTOajXDZVKw0xfebScKNVB7yuMOOG5CCYASBq
rCAPnmv7+eSgu7F9B+tw0yjEIsfmUKjTpe3IDTr3sPlryWnjBbJwqT8AvW1+5D0mtydLC/s3Y/R1
DGTC9l/ja5+KfXyaAqRi6B8kxrmSc5xGNjMhVsJMEXSzBbDksDmK5NmcClT/E46rJnP50X+6egZd
8zn+E+5+jNEg3OwHdDkOiNiDdyuV1AeeOkeQ6yDezck9FfMSl+JRwOyo/cQ0K+dChz9NyuBLrsWb
LLTVH+5vtbiDz0fSqoZTZjkTOCC1+HMAt9H3L6wslwjwdoKNXRYNRFTt99bztyGo8CESEynCRvN4
pBzLfthbd60rC8wTgsjhAbcEvmk9qZbNcwf6YP7W4jcEU8fUDdwVGVbNVCZUVn9Xze+rZG3usqGr
fptt7FA1g2VisgOMfkCvWsYWHE/1O8/DfO6URJfbRanru5t/lRUNEA0gC0WRA8t7uTt/c53vl0tN
u/xBk3eNgxhSkYfd1leqmUb4jeTvbGSSKgRMEZI2H1wGUCTnykK7JS5iqDBU3BGCwxP2S3v7Wrgx
hNEK3X0EGIdYe8keB9+BYGbQWS6tbotpOvLFhWms+5gVI21pRFjeUtzq2V065EwRKbUOw00R/Vn4
vKPlTDWe7VBqnU3iz+YUzN9azDJDzW8UEa5QR4e/HhlX+c7PUSURyK2fm7fRY2mE30h8r8dHL6BD
Ue0WUxr/JOHZp9/BwOSI1LdIQ41NlHhRh4AHlAN55T0QK19nVT7kfAQfjm64jnYY3F2IMU1KYj+H
LqYmovt8zoDUS93pIycuAf0nri3cUNIYFuiJxjEONXi1zfDxu7qYbO3U8vsRMSgnOt66x4ODqqHA
F12YzMjGXBwXLwFnBJrVe9IlZo4F3y2FFrXlmn8l6TCT3Azqxc2KUyt5z8CM72pHS1nxwiXmmYtp
f1zLfaxDQwDnArUv7vFZ7RurJgBQOsjEQAHpGob399VfT+W1r5ZiD32ikfry+t1MDJnHOtu3zVyb
27+X/mP8Wp0ReHhsM7pDMIcghcwECmC889OXfYtlEFETlnrLECEybRuC04zRCv0KPT/87fBhEAmW
VdOxy/OaaabsGpNdUSrMKBB4JlI5kGfJmG+9+WIu/1URI9moh/jXbrVy9n0tVZjgQrso0iFoAJIq
qB59BOnOnBaWrlx08n6QSiHRYRjjGLuD7881EAxqQDhazE68MJZzgJzo9wptpEZDaV6LqQbxspzx
YybEUJGG7upBwShcEf68MaGfxBKJXPicRuk+HOaQFLkvwGffyO52zGfbjZ8jzUgolEpfMX2OiKgE
ZoYODUTxwPZe/KVrO9SdNq4xZw2NViYEbzp58CQym/FbcAAT4S/LDB7hCeCqYITjt2MY99o3Kvjt
PQPhUGZvk8i3ezyUOlosByBGhNW5aVHNOhGs6zqjuJDpfgTlI9J6Fdl9a/AkdCRzynrNmAgKFSDD
7tqGLg0DO7zKsgKLcSCHLkvrZZfcE7PW8QZqLi40hH3Wdd6rC/qLOxEVZjWRdIFw8Ceg9/dR1ysq
NkBvbCQkyVnqLKISh6/WmR1/oE9G3xegDM48VQD/Qrf6jJVmBcyfy4XxMjHeJQTYka/cw/Q46CaS
XmJzFCwTvroPh7DAvNZnh4rO+R48FjapnAQb4G9KXG/Pi4+aSPq8Pd2s40C+cupzoYGw361mOcnD
NUttjzwMYouCpHwTj9MxVxitXJxJxZEPbSVUWfOblCjqQXyBuzEffi9ju3OH+88HlTR9+LSn2bzp
nbbG6l+tiAbs93Eh39qwAK19lOJrLIfhNeZtH+Eb8gj8HUQjJwqFKVKz6f25y62JyGJskZdEl4yy
gv7+kEQOQ4UzCm7aw8z+2m5qg62octOYqablOlkl+40Fzp+mh40buEcJpsLjknzLh7ko/zudrGyh
7ysfnmGJFWcWUNYwgCxPh5V4bNxpmltIex+dCMRjMCM5nF2folLc+LAUqFbE3NzRTyS8KapdbIUJ
Pl5QJkI0ikUPuScckir5mcZBYEI2D1j30J5r7oNxlf+BSMC/+7g+6Wz60GUoRtMcPTnyuxXNkrKj
BfL4XMOCA1ZmRTrOo9jfn2MH87u74OJMyo4TBYxct6TDMQ/54eJfzFbijxFJq2O/6JcEcfgF6UJS
5s5GZ3pFbazTZ9AkwmYMLwZ1ucEbISkLV08f4Cn5KV/AbHmt/XtNz4dwYQbe3pPzVvLSuO0hBEww
rD2LF7IkUqannv5CKhXIEdv3fis/FSUDvAFsoJhR40XH2g+KgosN9pimkOIUAZRKAilV/HltXuyt
7BAS36KH3i7WI17PPITtGT7CI34ndQiDmS+Oj4cP3nRw8sd+aacnHI0PV4+VGdaUvbfeNkcGBUF+
tOQDddlwW1fPBlV0eBX3zPn9L2P4bqQFdN+cBP6HGrT8y6mbogsLX5VCoYtywgncjhhv35a1c8pS
P6YesCKn/fYT0OIWzIUEuugiPpbVVRZ/vYLMUlo4ABleZ+iOqft3emGd4LeGqXVVQ0limn9L469f
QwTmk1Nux3EPk3Jvznr+biV6ogPdOElEgxjl4JSQt4fLU3c3BDZc9mhEND8ggyvUSCPIQfRFnH4j
N11qeiEx6cDavIhcaFClDJ4tTjp0s0nMnhA2InN8dcsBsGdj06GC1iIMXw7VIDKXdeSotxDceYbN
kB4QV/sqxA3TlBeSTKw5B2wQRrVV/HZszpx1RsFWvlwyKJ4l1m1u7A1CSzOhdCCC5u/SOZAUApT9
9NHVhUD5QLC+gtOVxcqmxmxWBSb9rQ6B4Q7PyFh2Y6pk1A2+svyp11DE0CL2AsY6fJipQeVW9bDx
qM6GzI3OPQpN7OA2BOKA/DEr4sAcUkIxO/7f2q5/UJsRCYpsn0UfV8z6pcDt+Wbv0pV2Yy9lx4V/
AC5d0LbPJVPWUTNuJLADaRwy4jAG8ePBgI9kSHZTDk6yrVGq1BrNmTqEuowulshQhVzTYQacokFw
aZXsmO5Yo5fcaUVr71iXysf8GHuCIH/0JsLcw4MRf0CPwkvu4egLELOZtY2xRezNJsFFA+VTuoD4
Zbvx7jKOuL/hh5NFXnmiIwh+nCN9agaIxsZfN386iP3EfYDklAU7bAJ5yndvE79YS42X9S/g49Vw
hYHKbqgSPTxXe/6PvYrjGh1VMJr0lwuqFpuSxM44P6iMb8rXoNhrgXSHxZATjnO4dL1uQrcKe8uY
x7/tIAAWFhG2Kdbx6N9IyfhXpRCNG2N8vWa55oHA6uDzoBPZKFvoGHpqk44RrZVy5Dj7HzwDWvVX
QnIgumikBpDGfR/cC4tUV24RCtMvFOWlVODvGupc9Dk+eoff0Ytg2ZyhBKath+ZTE99HhC3HyMxg
bpXJpvZglQJxKmjuhglxcDbGsYWjVwzVJkAmFxH6HEbKyVOIENW2F5gY/7fPj0h5PJs8VLoTc2T1
S7W1vfKSj1AuM7cK3rvp2PGHJNiob27vS50p9D/zJCBC2fpv6an5wOxvKeLvvXqOWC4BGYnygzbH
wvA2ZI4cikII2F5swmpe0qrbdU5U4Mh/DxFT4LRXf7w86SxgeN5d3J7Pr5t6nGd2q6gd5p8LV/0Z
b/5mlsDArzYl3lhFYa4osWwpzh4ZnX6j7W6Cdg6R+w0R8TEUjazBrkHv5Mi+ZFCImYNAxlPz7wJQ
Cz4VefYJVO+5hOGps99Jb5Je/LcNY77jwUvRRZt7I6DgNbWswxKQNdQDjuA3WwuDjDxgjk+lvLX0
aP5XLh4daUcR2zB15ZV0h9C45/ow/gTqc20IL845CO6ILfQ/vC1xJjua7nw+ZQ70bx68Op/GuOXE
kJsc653YPQpcobP6aNCEn2zl0VVEgq8nrfWyoD7FLTdHZH852HyodhhfBpjCsEFlS7fdKJe9mWoM
z3UNOsp9VgFgZazX9fuGs8k9gP4XKtHyfoR+w1x4l4OndFrFQXI1iXoAdvHSvez3vcApF1bBf12L
b2CMkRE0KQof5u5xhACs3LY+rnxpllqYCznf+QKo52EP4wyVM4TLYZWeYU7zoI1+ZUS4hLcs84UQ
LLD8mOUM3Xo4jkQIRwGKJ6GLzVhurgfDnHtQSyVT7WJmXBaMYA0k19ZY6Y+5NFVzX7zUNyb8ruCv
O+d99jgh3G3b5SJDMpQxkqhx8NvBEx2U0NespabgoaoDjrLXPZjqiKppnsYu2agoFHwCWwNbAVcS
+/dRC/I6shg4FQgT2rcUpjVnakcfON4QstYfeu7hqVe3QUPy/VyTtnxUz11/+tsW/zmnFdEF2jmT
7YAlN9rvOa0UH3cYCHrIs97bTU+sNqsLHg7XJ2agviL6uE+mFd+xeaNmN9T+xZQwsVFNo7Qy/3ww
q+itnsnXkMX769Nnoc2a9kCJRE25B0brf1u/3gb/6bYuqH1eS0kcWP+kf0fgtnugmeO0zmbxVpZF
AW8ju4kcAoX28GUqvsnhKUvLuj0Ji6al2vALjEj8XeJ9IOMSQagnV+jD9MX4PIZ5E8o2pqReTsHW
/RO4habUf6UdYyfU4J38yBkzbAm31AF7DYt0hLMW0ijCPAgmuzgN2o8uhITmTZm424UArpLr5z92
F0o8HA6bG2RvEx+43xRWMwE1Np+RZ13zjoCF/Ryp0zDndpzziI9tgOe0cBDbBSGCah1JyTV83Mz+
Oru6GEAIroNMVe/39M07wvE5n1SLa/yV8iUFgrjSmJZ4GzdDRv+1MNoowM3dNf+rtUMkWNNYV6WV
sjvKqv2nSw88ZZMcuusi0r+yuFuRDLbhinlbaXL1NQtSmedVU1dhxh/95ZNdmU7Uqauaerefm/qP
YcAIuvPDDhcve8pCP71YeDiEGXoI4OEQxgkHWwuVDLepaDzPuNml7fMiGcgcyPHLccKtkCDH4DTR
xOBVdeOxijiD0nTqz6FrkC6cExoD6pk+0bkwkO/YNM92fdqkYnlDf/SKpHP57ymsFXrIT17gYGwV
JtTHr/FdbeMnQlrjUXXZC+QDnV+bNm5QYbuxUo2qZqlunWokilqYnTz12j51JWQeW9Xu/c7bAz6+
FTbRIBtAc6NCuFtVt50+ZFo7IQLirtxrjT8/F9o+HsWhe/fgdoXu7OtE+so3awe3bvwkUz9J6aiE
U8HQn+3ejlRrFNdaqhp++iQPHVF3wac7cgDEA3L5FLWlXIAUHiSx/gRWiYafy2ptwNBr3Z5opZbW
jb4a18LfUgHpaoMOrIT9KnEMlSOr4ehG2birnTM1p5M2w03Z0gWHs51k/LaC9QqVu7a40nl/YDSx
4txCDg/1kGuLjwcRx5Ya/balhVTsg1TdM6NVe9QG4ZZ7QNclQ7961kOTFUikrb2YzEVceK7lkpak
5SeFxHQ+ZKIIr2s46O9oq25faCB9y+HNuyrkxtWK7+DlYuA11cI5U0lrfICjkExwKzrBqyv66SU8
gbmI8cDLvlad+kPa+Ef6PQBWF1Nr5WyqUmw4e3EpYErroaBBr3OjrLiYKt7m3Qdm8fFVwbMQtK/q
8WXRFUcUPXkJsVIGenMZAQ+bTphnEO7031jg/7O1M7L9ICtQ1aYEWLfYnK05wHiYgInf3PeyFBIK
39yRQMRJU31MsqX9hZI9tjVeLrIzNEnGKFA3sYObI3dQ/HDc5m2BJ0McP0ZaNomLgLTDKDfvJIbD
YQpIntkUISXHvs6oCmE2KHcP5KJOzAZQIJpWEz7xJmgx6CA50LEne+2CtKlDvbPjDlRZvbbOdkYz
QOnTXC2o+nnkrTuauOwqH3gADISxDsojbkXTEuNi9hhQlZvIPlzA/6At9+ANxinGt4ukEOrj1Vy2
WlOQhspu1ucYAxqXav3nBjY4BpC/k0TSSiijrsVEM0Q2DBFsJkvf0408NGZ16qIgS9gG8twI/X/s
59rRkeVXJixDvdRsDMxOkvwbI2hDNgo5r4/afKykCpA1bSXNDdVqBiDN29GYiYMakiOre88al9Vh
QwiaE0sllLUdpKxD8ChvANuGdtoXL3tbScuczyH8OYsCE27pB5dbfWrDYBtq1W/OHeivk1bFnwbW
saDHuWQtBr+G9ILwDND9YZ4r+li+tyrLZBwHmaCUYFOzyPnMZbg1E7ujLMKx2mLcJv82S5OuEW6C
Ra2gDneoNfveRw0Yy5TbBAqLYxVrZ0IrzYyywCJ0Hy+PEaTC3CvhXJoW5uc2QU7dwFof0rgjI8Hn
lrDPMZvH1cEBNKgdXwu5HGAiovC4hP7EtETIiET5oVjR45nby6OVb46TAjH3HOdHnd63wOo9uQNU
LJ4cF82xd+fetmCXdMb2IpLImRf7+2tqq2mXvPRElfAeOmmI6482ISFN60ysAeHdnxhgfmyztrZK
VIb/+esAo+Nny8u2zAL49LqGtBHRRhLVJfYPDwa1WVA/+XBSiTyxkxoDtppJQ3TH6YicoNk7amuf
IJrFmBcMsSSnwhEBLU3q0b7iPeB/+XTC1gGW6ZADBnoIxF9KqM5MASX+FhlVWMCBZ2tE77Dx7t5u
Hj2hTcnGH+lP/6uRlwtGPL08MCnS0bQcpj5Yzl1DlIsTBjDJMrm7aqDtC8Jsp3GIiS1RBheE9qMM
ApICIIu31Q7G/1L+27oSN6c5SmnkzOXTaDGOI7sZL5W2F6LIG+M8xl7ShWegocJu63GtTUOsVHEr
Q7iuStD3DFCB2leq9iKh4Pu6v4opvKw2eATiGO+XWreVXBADbR/UdtKBWIxFO5VaEJhw4Pt8B/ky
9Fy9IgPMqhq7NOwYJnz8mmrUhY5Y4JE4WNtgWY6QPArw/lwDsEa6U4qk+k/onwxsqgTpUoTRkqCA
GW1i732YBrxxOFd00akaXDci79UGm0HP3nsVqrgtdBtv4lNlBUl68VRK6MAMHFuX51/osKJM1zyr
DE1Fya1Q8YKgvza1tLStsW0lEbRi/sJ3zk4FN6s+cWBQm8koBU4RSTpHYJp0lxA8C8HDE/cvEThM
ukUK2B9GnulT4rJpJH1SGb34nmoDMAzMJtKzBFvlKJi4XFzXQLygN8vM0hWoTrAGA+/3jPNRgHKB
x+k9G6LZ6dvZv3cUzs3xB5s6j+Ll+EgIXFaJfO0elrvJPmW0Mnj31o3bduX24Qq+jjCeQXW/TGR3
X7E7J4Mv+8j/xgad6rE2iMkMvJUf4yzohEeP4OWGfcsXr9PEv21yU6GbmvQCN5C2Q3+wAISargJ8
dCrtWWJ/Z1yrxnVAyjeA+rObA86+ArhpGlzFjuDjqvRPDlbXddZotgWOv0nmXelhn/DDJ5K3lRuy
DVFo6cYVmKuIOEqk6lSihp57qN22t4Kti3y4v9WWK71gP4QjaCgywHFVreoxEWY76eiz1pN/LcMX
3B79vsbbX9T7Jgu3peGrN/fC4K3g8Pcgajeuggtp5iJ1QEGMWAq7O6NSrkVeCpWY0o+Z9bNL/qJk
+rVpy8UqEaVxnbWLoZJcNqHeLiJn0FLgzC8MaN4JUriTvw7qXpgGRvuJ8NhzvX2IDJgeDjpBaj5y
QkkxegpwUevi1docCCyDKJ/KUfuZ+a7naFivtPKiyebdxlq683EuthAdW29RaoQ1mk+utv+MUtWZ
e7+wkQSXStC8vSBgEAgHWlJW5f4dEYpEvoJiMZT3yMvY3fd2pgLAcaE59xQ8uZ5vknkCBtd7MWNK
JJt6DK28BuVfy1xtyrpgVSetH1uI0z2VkxLTkodwcYwoVzcy8Si5iyPUhi2u7CGGGtSMQDLAJv/m
PpGWqt3pvZZi6Sn4wTIGRxJLqXlQfBxn42MJ1fUBVfQnxE+TfKpxuY4HceEeKbw1u0QK9WobIzHd
cPD9UlD6pq7JxeCJUm55duM30y2R8Dwf/JW/dL46zAcxmG9EcoLFFA0pE2gSJ/EfjozOpIfHnW0Z
H9Mi5E3szI7jYeP5jeCnccfjwPb/ZJkRI0c8UbEmPT2/PnW+fpGOv46bmMuZi3nPDEYaF4ssy7vg
Lc+57d7tBub3P0+WkcmrG/ZegmW0vsoG1GqUBa4e+p2iAwLqghGiWCbQ1Wv1Q0ditWeW6tVjdVls
1oRizYVwHx80j3VvQjV+jeMMRoEXrZbNhPC3wmpd52Y6cnLmhY8vWToBH92vLjxMrJciEzViDD3Y
KgvS8nP8/D28j9StoHaAFGFSC5Hn3QhUjJypWdT5uf+krKV5H2DBCvbI9zni3J8Oh5Q9/JBLUE6s
PqF/+0Q7g6+Uq/DAt7X4rjKagCxH0Hj7FfiA635Fil0JdCb2/v4AASKztEjo+5FtLutOWyQZxilz
Mop6SfEC+9LSlVlgV616L0lS6+orW5ecscM4/YjPKuE1v9XkDniabFzv60ZqxezkOR8LpNvzcbDX
7BAxRFsRkDhg8ioE8nqXnOWtqqL5onOtZj0wjwMJn/r+mc+9qf6GsCaxNqeV0Qfb0NFV76QxpZjP
joJk8NmotNAsQG/Liwkirxw4wudqA11kjJKWLJ/1VkxU5Zkv8mz5z5chgItA5xnqrT/AjfGr2A2Z
vpIl3SCDTwb9jbYdNbEn017RzaCEaBPMoCW6gD4jwMAdOpEIYiZuofmEZjjE1HGYS0UUTHMKmexu
IDntqCXoJQUWj92CLQ7XsadG4JvwjzupbZ0pNaKQjJiwGStsby19KlqxVrzwC8jnQMINot07/FQV
ngN5xE0LWOFIuG7Dw48BBMPj7ZtPwpGsEaZH79lpyACiTfUP6cCchZ/6dOM75sUAxC0Bob5O+Qg7
KXFmrz97Vg7xOEzfGnwrQeZ/3ExZwdLoS0/u9hyuZvalNo9rhe2IMGhGIEC1lWe0+Pa1HCDBHOXb
KDrJc4MSxwBbjq+VIBgUmh7WvB1A8Fa5TrETKMp7Ksm0bNWxjC5sADVrQ8/eL5TY+jFCiM71usQk
3dPIP8WccslO6/uTZORtoFTJ5rQq09Xp38YfBSDTCAkOHmIdcuht/PWrRkf15tefDt0tkTj/GIvx
73a56AZeoNFe//9hidh8JFUTdY7QvuZ4doYJpMEYaR6UXVpKnPa9Uf8RybiGPzhBl8l5i9cFMxBG
23jD5lFNIDha1NiUo1AP+5OEb1i6BB1t7Ne8SJ6ghqW6B/fG9r0iAMPqb8GZtqMGCp3o3K+mQqMJ
5Ii5wtbyNE9ycbh7mkiIoQL7i0vmivVnA6ajz710P1bKhhVq5GwOz080aYn5EF7CoVg90KH2Lolq
UJ3a6ruos/Fbi5FzSIMt0zktdQnL0XGjTpnK7YHLUH+BebPkiUt/PFIo5xcsneX+4yNW6fqbw2H6
C2VHYr7MFwmRz25d+x1CjrPYSqaPGfqK2hZxxbnlnlbG5xwrz8wM/V2enWloUDYWMSu9k6styecg
fdArBD8oBevdqu7d9Sg93aM5FgxJtQRg55+dXf5xIiqNwNtJ/QBIAZPGUwPDcD3rO78L1e7plLbK
/Eor013DFg6HjZpUV/FgjkdPpSkC9bKBiDUmjRlWU+TlHYnWAn9TfM2fCLGBFg/NOJgD2iogxPlv
GNVeBqNwb0mSl332u5Jia8kuM0afA5dVPLYmu2NoH3wB40ZBs6QiP9Rsm6INLS3Dt4LZr7DKnu1x
Y1CFrxHdAdMa+BpnuJ6JW5PfHyLGrmqS0e9uG9vxm+30dEna4R6V0EL/gYyt6dfMkKrkgrRTFd90
4TjXcQH1EyQxfNrFWgRBGMwI1hBEylGZF+ZRnHbmAfMbb2aPO+pSNNPeAHmAcFqWzAqiE6YqaHdS
9/mGbihnenpw4dx0VvwNTJttF1tloMSD+YgkCdyXJttepGGYf9cJ/Ogv+JK2py+mrE1j6zjSZh3w
jgvnyQZMHh1LPSGReSl5RaNvLqBAjycVlmPvSFWlimw5Z1t3CI/hlxB11UphVkJzuWi2umwQwe7K
Diu/t4uVNcRWIWlQN2C/kW5il/gDnfMoKrdToGwsobt26GuyZv4t9CsUM8QUash8WnW1F528u6HJ
3uc4TT2H/abYA0efPFCW+JHvXSXCxV9tlGQ4MSMY9MR04kZi1hk612VVHmApdEWGW3WNprrCDSop
FG0D95aMHSMct94xjjm0NjVQr7Qil/JGJiSv7JLXDUcuwskKOWyt2hxuv1UTevzh1rXsyG/hvVYh
90j3xDL/28itg9CXmkPYninowdmmi0kob+Jmuq+m8QsTYFO9MO1aY3AuMsuAjERiL68Avsnqbc/v
zR39CBLq0seQBR2ic2kdhsMWbq0OpfQOOvoHq6oN2BFw8Ohp1SF0kVfzkhMM6RXLRKxR92/3m4cq
EWCsFXPrsxgPYNQp2xDDcW2eGowUQ1U/yEdH8rLmrx9/xiFq1oqJB/LZmMkfgmwvFCP/zUSbQ8Cy
29bwyvZoeiFprGJUWqNTIxgP7KCOu7ABxv5CuuYQx5ipQq4xb5VqIEjy8ZyicvOWL/KfO9ZaFE1L
1lMKAxR7WOnyEwpRHRUINlNyMrYcBGw5Bka1Wg7BONWHf7quPp86WR1mg+MvUamNZ/kaV8yyC8iW
fB0t5FSWOFbLbPK0UEs7sK/L2A1k+I/gZ9yamX+IjHkotWZGIw2142CG1cEVHwHKlL3/81/MtYRy
kseCYUel9wXdbi5E12N/9AHlyeirs2/nSaHuSCIwf3xM2vzIyfIcjPbBjFKkBhIw8PIvEtgllSoD
YAZGJJa/EiOfRdp5sgnx27NOceLVrYRMN91JiVo56E3lTukVmHfd6aWet+lku66JKiKsErqWrj/9
NLMKQ5TNpVoxGHj1Tcm5F4hUylLfuIGkMrMpFFxboqtIt27+gbbNBcN+eCSwzc71Vx/gM18j4Rc5
BWynwFutA/wvy2rNHBV4XsUtc/KNic+ZVL3RJ3tSZva7bR93aOpTC2nzJR13xuQBDNxLTPubdhPa
gtL+IMiM5l0aHFiUXjh3iBVdAiJFeYqzrF4nYmCgJS7+AjHUrsDhQ4X/+MqZY3RGKQ8CFub+Isnm
Lgs+6SS8RK+MthgT9qZ3X0CWJ/UOWAgKsMBqn1YCbyp7OrFryv0uslGVnvcqErBU1P2xUn+uWiUj
ib7BTU09E2VJnuRsXaG+ZKgwBNbKjUFcL6mV34dw9p5qs4haMxk6HiettXpP4SaKJH4SYq9+DNZ0
liqHCbZYSE+Y7AqbTqeR+fE7EmOpu6MYNUmsgxHj30uQm1v0juFZKezRA2Ado7KRYD4ONddJ+3Kh
uL/mkhr1ECpUZi1NOSsovR0pOJ2QRz7olnPlPKe3juowtwhSsnWuFxxEHZGSXQMbxr5o2Cx7KABN
Iutr/sF7z2Ftb0G/qcCYA49k3qtLEkq/CLd1DWFu+j/Kg+AD/7K5z/A1+W6/Rgoh3RYjXerawGPV
jF2QX/5GjAfq7jYlmvmQ/PUFSdrKGgXqbKNKMFKPIeKEtEKNgyUZmoyLGEQemic6UdxQi4cL0nJz
M1TfqsuZjlFK/yfPE9LW1Tt4mkEiH3gCrRpDG3S+AvXtkWC2EAwCJAEueHeDrk5aTFrl1n6X6lC3
wFtvpDRDyyWfKq5l8uwYTuuXvxVvKgusNBlbWTrXjo+BYSq3kGA8cxJfAr74156sbWkjLKHwXyDM
QgpPDSIeS/0lYqguNX3R18hYWwljjvWsBqE+K5Z40o1ycNr2zwoFc7izqL11UARw+dyggddkmrLX
8LS9cM9rl7AyqKxxIR0u4bZi5Hg41uYShXrqyWtRtFHqmruMPcoJLWhLim8lPG4K3dn76oXI6nhX
EgOyekhqLtdtEsLRiNntsBBCJ/dV0TDiN2w45mzlMr4d9r93ocHSaHfdx0yW2ByPmMuuV36oTRGY
Lpwma08ceRYsgcMbeptOAQbO2GtqN7zwe5JKRxeAkA0/UDS59EZ72ZIY5OCNiap7R53ebjYQLXq9
1Oq0Kv/UBLpLZLT8KP1d/zf7QL3W/ycxGIYbEu+2dd+CQHueiXVSPPZF6h8ylZMEob7sgtcAejO1
mOvlzAfs0uAQZ5kxhAPB+Na2zR8yugBUaJA5rTRRHY1eFCTZx9TvaWxexKM0gvHNCHOBpXnrNpzz
dgZRgU5B3xszpiIiwl1A55PpSqdAEmO5vBb7JZ+1jQY0BumHe7h9brz+EvjUBo8LH2oFb7zWnS0i
RsuUMW4Ywo6W03XYr2wkvf4tTom8lxb7/YzPGrAqD6QFIv3CbPWgNuSWVSDxToDQhMnxW8d2rB52
cy2Ej73LOt6MtBFudC1dYD+WoxaIv2UOGmuWX1CZEFRIda1ii7RDqWfaVOTW+dj2E3o5XgQqPU0G
tBNj/PyQVzTkLFWIwcTOIeYWsplH8U/3opKK0BUPBSMm7a1QiH8c5/s7ygqqQuCLdZQBKNifAS6k
DO3IVWYO0L2IMVOb3GeL1X9gqcwuoZHoc2HsaMkcdeH3FWI8/s1Swi4vdy+/QY1xQuVaG9iptzlm
6vyLeFzDrkHHL/NW7Mp+nqWzgBG8MyK+5AaVMNtgfRY1uygKwWp2q6o8q6EjlSDfwPKH8f/TSvdS
3t+ihCOKUz8gklm1euDBMUO+6Q5BObFPbxQw1qhxsbzP8heW0C8HzjGfztnvoXs3n6GBarz5C2Ve
sGeaNvAwf4V7QXC2udPCLR/8SjdaU5pYyFaJ3N202U98D7vLhfbnd0V9i2h4cWzN6oaIOj37IDv2
EMF3yySiyEwLTBnp9aD3PtlKmfFj2SAFuE7Lu43hYdGSEZjsNzd46ujH5y0rUZCcQAT6AF/AifPQ
o6sUZpdt1A4W4i6S90UpUwR6qPXfvQt6jFFcn550Nkp9Zu92EDExiXiFq2L5JNi9rxbdARUZlU7s
w3qQP05oDIIacA9FBh5oc9C1ZraZPfqrmzp7vjMqBR9OLjXfj+ay98IgGuoeh5SQ/z44WdT3VQ7G
ABKuVvg+/5wIFtWS7X2n5oS6kcgFfB2P12/EE9ifYDWEd8+moJGxVIyk7z2tQLXPDryVD8dH8CDM
y+EJbIY2rzHQ7nD9/kzChRweEz5CnIt+fmgG8j4u+2qnGgjZv4zPjh6x650PrOg28vSlv+r2/8DZ
kLcZ1WZahOLQHi3jBQwjmS5/oInVxobtgWsZmmoN5rF43R/YeQ0LrfBVwZbbh+3FEDRMlVi7V5AU
GRgC0mY4CyTKC8b/ZDm5qBDnyE/YeEV1L56H83kifCareAcBCiD2bu92WkLTQh+YKBmw2LlT7gyf
eEgoO46Gn9FgBFl2FpTeDfKam9KcCJSesFOllGzfZ/soEpHyPOwJBOek7+JEDpta+ghU6oOvcJa2
BWAlPkl9ScPH6wLeC2A5WC9eVkxRqOSUA3F/fz4NfFPWvnzJfnDj8oWyDLjsXkz23dKGZWF1OFEi
kVswqE0bMm6dTQVhRmmdG5K0UJPsIG2IPSp8flYIMzCCP7aCRvpU3n83nraOIWVHYSvtNKiGGyZB
ashiUhsus99nRzCfa/ZDH/kYkrVA4h1rZN1ZRQz0HjIRyoGMTRqHGxR3JlCRuNFEbChF1wxPO+gc
r9wuz8Kqn87QEE0jJvv/v8sbYxNBrivNQ93xB0Cm3yqlh5FBJPyMK+CgugLeOxavk2h0FLZBOFsY
UzwePTaySUxksnNPypzWY/jPRBn/Cv5t890IO40ONskZYnAlpnnBQVGr2RvaFqq+WQx54bmPsaYv
3Qay7MpuNxPGalbvyaXxJCSO1OBpybsQonArsDm9Ku4mvEYdU6+XHA7t+n8lfptoyGupn6X2rwsf
4EiHHX1qp8zyFKJ4aaUxc5aDy+pMkHWxjsZR7CpLyCqak/uPHXZEBvaXXws5eKejUkIH/4/ai3P4
cY05CjEdFN6qXhE7C16mVp2W3ZvfCiL1Dqw+UYAnw+dQ2FoyXfiMSshDu0P2A81U22sKvSD4GfNc
7VAS5KE2iAGPFyw3WiJaHuqXEPl3nEyUMceGJkL37WJXDfNGfYVc3jextYTvPj2IfAJfm/1QU5jQ
ugTfG6bfOJcx+3c0stM6zdWBUX7rBi87BPx9nPcvXb+TWJWHcgY5+iZD1I3bTOoN0mZ2NIZN6mXU
jfyrrk3wXNsROl8HfY8extJD1sOBAQwvsifz0VHl+JnJFB7qJODGob3CQ5r2S9uAvEk3rHRxA+EV
sH9I8vUee1ElDGRKV9h3/XMeT1UU5vspn0QVpKf6mL72Yv05sdeu8oCOldjiSJLg/wpN75murntF
4fxwO/TRhQziifkX4YwPTOcyg3OZsFbKMOY56gW+ZY/fJVc+GXTlzA5nRCSieIiagS1d9nZ8P4u7
dTv5pUQMN3lc+n2JkR3HN34pnxs5WH9bAVXLvtFTpPV/yvMLurEkgSGOdc1TVpFra023MyYzQ0Jf
p6dc/0Xa0wuo16/i/EMQTnTDkIi+FiI7n26V5gLFiBdLL+evhuSkRLrw363RCZcQ2+zlHXCBZcea
sU9HEXmZcmB9tKBYm2O615I4QrF+rX18XQrlWfks7H4Q/6qI/CjM++0kcC+dl7LiQw6TKOEqFhCK
x9ORGVv1HvnqeKNjYGcon6bGI86Otha5EAQJe4jGI7OvIeAWgoGIHGZsKQpd4QFKRnlw8zE5BAho
kq84vVDxbVE7yrDGirX7dH6Fs6ikyKga2q9xDW0KL5Sa8HEiKnq9xI99lplSJTFCJAerSiW7gROy
KwnSbRQ2VQp6PJpe0BIykZVKAY9Marf56SR425enhD/5crwvV2ay4gEJmNCLIz0f2/ZBhq1ZvVuO
xVw9mEDaHpAQsKyKWup2THpX7Agx5a/nLfxzh+I0zbkEjUO2nhpsWuGPdHr+hi3m5pRKZrpaXc6u
2XFnwfxFYwjNBOCKEKxzLhWrXU6ejZEQHeNyPKcOzMY32hPV8QdI7+54AuQwwWFJXGSrDMAWR9Su
so1jBId2FE4+eecxohYryWqRio70FLtCe/XpZuY8lqN0Cbn45RJzAkRUUB7kb5b0Qafk8pag9J+O
RZqMEVJb4kNdEQeOT4jfCc4WK0rvR/0PjMoWdr/u9+HMeualUC61EzT6+Fd8bMx1bp2MQwH9FKyh
zW8y22rGwKqc32SuZZ8+53iUqkB53z2t7dgVQmdJxLE/uguVrQP4xw1qA5cHDQc518xAubeGP39X
7BJi7lIqUnJQ/bgveRlQ9t/fxlEypg7LMHjCl573LxA9NAQNTpybY65Pan+CIFBxp//b1ctL0w7/
hWLHyVsALq42SRZBbJSB+WQvXGn1Ww7RWelpRjOp1YBdiIBQoPMeW+ws8nCVOiqM5rVWa0/mcDa9
7a1L+B/Wn/cXBiix1nzC2vkhZqIOyTge+jvnLJO7t3x6kcNvtwN58YqeRDeP+VpX8K9mprTFde8j
W2KnnMfvBQyM5YmaGF+WaXLJ7LvMTtGJXf3E/VXGyf7pwLVRBIcdcWTqfAEZl6hUohtWXz7+YLup
HX6E2eyflGsVeVxqPBGsGUTibAnspJT9zAbsyt2537G22mau4YJBvdHvI8+PfImQzk/Uui6rGKvZ
iKY21J2GQakufiKafW9nLCpo8UW+qt8IfZp1yMUGQXt+px/KqQIwMHCl7CHmVRP9ERvRAVH7imKK
JSi7XfgvnIrZM5FLtVoEfTOuXxByNUryU0mYEYUkw+Nisq3KIHPYOE5alZvymdE0CF6LSfN0Bp/c
Wr1ye242ls0eWaauz6UCgoXlg/M0Beb0qdkbOrvkO1v/iCNfGpKLAnmW+QpuffIykgsDlLMKqKFN
9QANkaOpaFw/p3rIBeFnaEYKdrNhbYvzLoONzA/xo/WDVqNQQtSFHnMgLHOvwvq9tcewA/k6lHRB
4enMIlVQQCG2m1FjVfeQ4dlotPOLdtIuAEKv7uXWzlPC9y4JKoh6lHK21GsrY27st0GP4STeUjLL
N5KmZ49Z1yep1eJqdqnLaYcZo1qXFFMjGGEQHEH2z3kJRPbWLvtGi0hwgLeqWCLfTsAkzmMnLRlN
ojT8s8VuhiRwScg8xnxbe1HcOdBIfVLbsOAfQAkrvWeLoLEH3Xhy3aZbbEiPtCtB5koK/+R75t36
Au7Ne1zxwlb6WCoMJwyFgrYv1BMWa1NEOz86+nykLzqA3SWX4AlnjAtXlG5DEpXNmTP9jA6hM6/E
rBS6t4Jsb6PqOQchBH/ZJEEUXWrB0vttb8CIctREdkKge1b88BnuapDItAY9WepGXJeEUPzPGq6N
sM0dZCEq30o9OxC3Blpw/eIhLfp3fwqrwnl9Vm7QVR/pQQqIDRNeNHIq2lWPhRnvd0APiVgV91mN
YUTB5n3Mm89qCE6ckQ9vHN7QmJbJrg/eP+9URcMKH820NIwXBNl74fyprLW1byaOr7XAIOAI18Hn
eQ0sVAWLjK9H+wJsvR80NTxdKMVBYj2Kz0mGdlUtErbWHoRcbRriVmyEO1FveHVFqf42MsPM7PFB
cUHaiHufN71NQeezeR66z6gaZrUF4wHcJJZIC1eYOGAN9MA55dxRqRDe1UDmFBv4NARdIBnETk91
wptxsVHv8Sv+NoLuuVKuVpOSTOcpgNp7XRmj2Kf9nR+rGBz1zUcsPdAfBXRFMJIHc17aXgzaSkAL
9CNYKxGCJcVt0UGaYOaiPpAfpNdH3VCkIhAa2oSDfbIf4SZgXew/h+XTmF3T6xaLxdyTy368RTWq
w4tQ85XfFsiJ+K7DOt/XUPQHtDGEUaXVsBBifdMz53eZdiP9+54n3Pf17WMi1llvzU4CBcvJDOym
HuT0wHKYNsAMilvkiJlO74HmE4fW9j7XOaPNW05LEKnvMyka0h273naY0nCwxzLik/vI8+cX1BA5
5KSOBgIRn+Bs1lysjE0cc0V0bcB8jtin1DB9752VCoOKpcdGeRChirmJt1bjST8Rc1P3juEKq/xt
i3q7LUWMIDxJvnoeV24GtA1ctYDkwmS70kCkUrx+I6fgXVsQnxsCJrAPZcU4P6ebXabvWip/sgGA
+w/d1n/AxM6gE9wkRIo0T0rBspI44JriJcXNoYzI4hS1159hsfnTWIyyidQZ4Ue0olMq7OroAgAG
xOBseZk1zN28H2rt1c7UgIXZ/uQLWHcDJ8raWduDSqTzM2xZLfOI+v8MSt8vQCMkmNQcFrozG3S0
r7uBmw8f5iLy8XWRLaI92lIsUk/feYMB6qbjKr7PVVs+5HMdjKoJXklEtYJPJ8eyYZvzLxuGq6ar
68jUeI/de94jaKiTynzlZm2eqT67dgVk51+dhzlOByhvKhJD5s79i6SIjLMUwucqm0MBRnWSMcyn
aBmsRCBHkAoIpD/KbaRJL8l8Bx9AaUUtKD+ws55jRGU/7I3iTlahgTY2A7qItYU1hiFwCUIKvQlL
BqeJj7ZVaSP8uM6Ip3OjpquiNyi+XY0F5JDhdsOHq4qQf50PvKG6KqYnfOuOMBaA2SbsbOpFCnUB
USU/WiwJX6QB1pQF5MzZA9o0tDIYsKCfR4oIJoZTQiQ4h5v1CFRDrlndjyEkST3UpQ5A0BRsLeDx
QabkeriKokjW99S60XY5RWQMzRhcfriiFRNbay8Q8C+dNdRqqb8TgQ3SyZfEVtP0YXXEg56m3oyH
iTt1oNqtDwYGRc9sc0YSoJbt13WVuCiZv+2McTR/oIj8iJwo8MH+QhcGqtdsIZo15ZgrGA/DRaUi
pxRr2rtHphiIivSTn8iSrRh9nTVqoU8302GDsS3Mcjt8X81fXqjdxQ7+pUWP+HThNW2RvoMNwCLZ
LlUmmJWVgcQwJtdFZY66Fcyrli4VmnK58ezm2ssak2p0f8mj3NajhGg3epLNWgYAKqEAmu2mvB3w
iYhv2cU0t+VZah0P7Bv05a2tDn270YMIuUcQIRxh2meUfl5a4CeFkb0SbuEEsPpZ69lMFHynhc4M
1KJLi0Qg5AelLkeYb9gVWa6YxBh6jNtuSqVIy1N0OR1fsrQE2NtOIsfM12oDNxLcb2tHuUXD6ZLd
rW165f0pwtZmMkxglItx5DuSjUAFBEhIdy4RL6WJyM5Qehuj9dc8JZ28RSkkuq93xOJfFsEBsFQg
Z87Rpc2srXf60O5j9ZCTAgMd5Anvv2aRW8d/J/PxX0G3drTXndXY4SbdDUTSqd+cKig0jT9OJ4jk
kArrxLigznGfPliQw0ULX2/ZPgf/vbI+zoTA4xEXhaUoKTjfgpTlxlzsSgdb/IMC0U2slnA1LIye
3NH7Zrd3HdSI+ZZC8i94iSakr0okMfyXo4Ab/4pkdp66MDqPYRnKyLxaa/rGl0nB+YOtPQrg0GGM
FVEtfjBzCaoRFSoUHVkbJPSB7je9865ct/Phm1dQvqCSENB8GtwlHpJp350ja9/PrpA80qPJmOyO
psqBSUWFsVkKkFPw0bs0uTFmwzz/nU1gybzlCkEQ2lJjg/pStBhFmoEBU7kv53pzk23GU2DAl/Qv
nibZX5EucD/XuZnBO/Epur25IhyDtXJY9MaSWUHjc6M7EBaVE4TAvmo2o5SUE6TysVZAKhVEoF9L
an5KE0CchyuKFjPW6KxIiP6Z2WFNyMuLeMVAqwYicDoxKGEXY7s4mfAlkj23feORkjnsxXNP/+F+
crLHDnhzrom7myjBdMlkISvDYn2Nm564/uMg3c/Pl6hMloNMr0ReWrgYDfLKDSoeV2Rdz1m4qlUB
CcVw4ie0dmxF0ceesd7j5ogKvEZMITeDY6DG5x2/28UhNNTojHZN86LBGksW4FCBGh8CW/sV3bOV
wQ9mO0TiLfYuPsuokGsQf2NQzWlVmIMHzFJW9MkgSbLJLkkGYYJq2zPqmysnDFp6Fy8Z86b2x7RO
YsSrTUHhp8yrg/QlX1HBk0jtz3Dpt1JWhkAAVs2kUJhuetAScXJm8A/ZE9PJdhSbdZksIjvXqUl4
A9cNhMcn6DheSxnx1bNT6jumgAkuq98xEh9AL++WxnWQ714RZfjUAwErX+w1FeL7ovwrMwRHutXS
/V6l761FGKoNJccBvsm4oKC7yrmQ0iIBCcYKt3Bxn91iuPca1Z+7AAU1Vnu+cmkCxMXc2vUX5PiY
h+aXOAD3NJ/2b421d4Bxerrb8uIPcdF4NaEtmGoBBSCMymp9vEPc7WikKSs42Oz0kCNOMJfzVz4T
3G/EnPQHPT4PMvzhUC3VrdF1i4ZE28cyjP077IZvWRUkUZmJbSHoqkLY5kJBBGvzLPKwJn01KfUu
t1LDlO9wvZgN9Dk56OxmNQbo9oLJWPo6NFQL1bc/I7G2PXCl+CZv1hxoD+RYpjHi+rC1AARiKEUu
iNJm1EW/5jQK4xlxInqmfikJtlgJnKtS/RuP0167fyBeBWDqjlnr7D61FrpDo4L16J+Vgrz8bASP
haoDahEG8O+xR/6Y0jp0THIaT0637qSzV73ZoU0PGVcUtSdX2012n5a91/BLDe4W7qTpfdy48kz1
zgJL7hhXTx+wzucpUv5Mwaf+28nzsiYAfTOLVDdkTyhR4Ua8L6kD7c6JXwai1L7FlDyhHd/QsO5d
WZjLxXcWz39iOWColV3c/BhalRhjoe2tEoKMnqVxzKgXGRoXhkwBNHOK6wEEKotgF1hh6s3ECbMd
Bgf9SV6UkQaaYLWAhShEHM0E9AKtu9+MU4waMnE/wt+doe5D+jhC7QO1FShBfSJwaPx3IYDSiwaY
iGdLSeHrNAGWl9b1aRsrrLnv6iHVxGNUjBdYdxwwqMRdDBkNiPR9RfItEicWiTJDYFWaD/3tXRUp
89lvygzhryBGSCeSLTHS63kkW5WC2BrMWRHq3emphjAob0IRNeef5/67uwCLUVlDYhfvLrplXO5e
cOrPyxz04lArQujO7kxXit7u1DruTLYdC+Ta2cuLzq6uaLpHnwebPEvZi2ooMunqoUzfLExDRmtA
cJxosrgOllup7qPsFEdm/mpfc76vDnPAvAaslbqFI1UE0RIEcpzNiPIbIO99GOTG7lBLa3RsFREz
/ZIfgLhzAz9agCqyXJxqTwoNJkrd9HJ6ISekDOnQDojm1wyR4+bn1O5IM3KfPO8lWRfl5+FwE8TH
6o00C+pWB6tPnRZzQneb4mkoMwdZK2BPIdCXCnEWsOUiN1mMznMB6VO4O9EPyoy+GdlGkYW4hfGw
agNZqvVfuwn2tqLYUdFVKK1yhpcXDdDEUobNpfU094Hc9ARE9cp7uFIk539BpRm0buhjJZZPEWTN
54iDRTowCWowoe9hFfJ7kQ6KCey5AwcnPJfAbr9wmT11Kzoh7eNhIZJcto7QmiEcKdzm3kSpTyRF
J3bBxlHu8i//eeX2e4D0DqCiXscvJPUt7zfJWODa/sOElPMT1801AY7eNR3A2Tqn5ol6HfuIkJYa
6rRZryQGqp4rWTb7dAgF8joRvI+jI64oT8mEjViTbcj0DcC/2/kLwlQyhrA+x2S04kMclgvbq6ds
qpetsC4l5+iHmbzCM1Du9Z2pkPJaX1KcAuxkvVRzUHpgmLWaGNrtDjQAPnoslH+8bBx/bMkYHRfx
zgNUZHeyF83jnS7U+4ZtBtKpb1K2P5xfT7EnOdozBtgafPJcp0Bp9FrqQGjq6rUX4wSFNi5VAcCe
JO35VZUuF4KvgbaIJ+fdiFBCwGTVV2EyDODOo8MKgTJKMBHvKdkuzyzACCLnTLGKbndlKzX5mD/4
xuMEYGH9SEvvnapUEGRFUM3VfnAuMSMIsPNvfiCtFAY3W6hWFtLqUvY0H+4/4y5l9sm09KfPjg+/
0XPRDVMTDXkbS2slDluoNoU53bfhEweECmWK/dFWDetU4wzVQH92NCyJmE24eoLGdJAztdFk4nAS
6K6NtljJNdo0YpwpAIUgYpeWKRmLUUfqtTR5k4eJlbAZC3WG24X3dfE4PTFbiHKCLUkAv9xSI5tw
kbWGRRWaQHAkU0xORGQqEo4YdZ5KQoxZhDfdKQQjEIrraMdTeMxkhtwFrN6YgTsusNJ3EQxq7IXX
RM6lWmEYQBzhKj0d8/b/NTtOPQSxOKaxmNUGAVioN0FIZBdmUQe0EfQYcLk/P2EetwpctAUgx/eR
0Uy++ogUK2RTsBGc/hf4FGRIydmqqZ23jyKW1zsBw34z7HM28hfwEVoC4QCwPNvhfKAVmuPVDqgo
OHZ6gmUZYEAURn0F+L0qRu4bBErcySnDzQcnKYL6xKR0Cvl++OlPH/xWTkJ4Rd86JqeGvWorLYt+
YCGpZcy0bUUsQX2Q2/aXoQeUUXIQNvs6z42fOO4S4muT9kFNdLjyDUVMS7Kl3wJxjmO+fYujbhMs
x2bHtgFuoU58m/jIsNzGzTEMOAtc5Irpk+i7jiYtKRG9nzDShEiLXZnQx6kISEvT9Z6HuuAjnXJa
3xdKYt0FgevLot7wIwuJUeAEmYGvjNyrdGD2NV/leWzagEixNVdVqWgDbTOcmlF0LKZHd8awoot6
I+uiy6YmoT4HtM7u2hUSRflZpLM+hekr1m7CJFXXmhDeyxt0uMHQVz1Kv4YIZwKfCN/vZpGtu6AW
bTcDw1KMMGOkIbEXSbR9VgdnCeI1tqgcaF32KfwkaAkYnJL5EV02UpCi8Y0XdMt0tlYAQ00tWwi0
SqxE6HKUVljUyLesGSmgrX8irMwKMZQSsOPmFY6cca9B0CrAM2hvJiBogYTwqomfToknFloo7ZlH
DZQ5EAzFe+WEaFeNZa4NPrwxwqwWH0QWWcIQXhzTxWvLy7bF5mbjshw/qkKj5Sl1MC5kZN2eMn/U
fB/NeUyesHGaPddNlvW5HwA5t6eUneiK0EmF4Kgj1DM4Lt04hKT7kykHRhEPj10C23Ca1muEec0S
eox2Lhvpx63ZMCdLWif2eNc7dPe3eEWdjIEaQj5nAPldnLcOgeSfXp2AnjLbWQGagm/M9U8TtGgZ
Hub4FKlecHdlsoRnSopzfpNgNVDgjZ0iY7XVkwVDYrPvI8zoyzctLI46PPhD73nIioilgp3x910p
bIfzaCbu49KovXFiReWsYcQirJQb+SrkmQm7boUNzXP61LOZeU/TNBXQRrsd8UFxjSn5Ys6Dl2Cw
ZJE9F3BBoeIFLWarZXlj5zyMKE4I/E5WHBQBDOsEGiyzmIbZkuybHqGZX+XhP5OX4C54Dwh1bWkr
s9bSVKjuoizmXQ81HbzYgTjuj4YRLzbufPGzYa0oYa+vj3h/3jF8+aVIeybcjcVaYqI0mqAgxFg8
ATIriYZEjw4GRaL6qJBCTSqw6F3d2bZm26fRYYWdddlsfRg6fF9Fak4/h9fL1+4ZA5WQMi60YKrt
nuZXq8eE+LbKEw8dHqs/5RtBPwvCD7hIDopQ1JKQrSAaepn/R3GC4dLBTFDQEspnS4OWSrNJ6nrE
/l7cEgfzFZmrtPueaDMxNXDzmb0m33cbr2QDcKdhC/T6tKqdGt+WglqOAPBE/3Ruoz5lsZX8Mjbq
K2F1YTZYD3v1cITpxNFc1KcKoARXnghLvMrNQa5UeNj950sPXjLvoVhacfU41PJdhgis6cLfX42f
ThqcVs/OocsB9Q1HOquk0EhcT/aYgGaAj58BtLtLGWPBmJNrMvxLlapkPA+GIEJu69xfaDHEgcel
4iqBycTgHYi7HA2OeO10A+tDscZJWm6H7e2li6GiCAiKC7S19gSytF25ntxgOVTfDWQpYTbZGMA3
++ZI1WclLGHi+UlRt+9aWRPzDJevpvZqi3h3mzRnw4Q1ITSvSSMufql6PNOrft81kN/Qv1FbB63K
5UPXDXb/gMcGxYHO4iQ+0XBqfltMxsPDAzp60nuQBFC4ksCyiHiApw2gEJ5Eb4RywM4Ps8Zu9EtM
A4im375GrMltqS/l0in9GIsc2m4R80tEsMhhdEG5MbsTAVoMxi6PbPmXff0VeFiLgJni4CWxdSbf
l7Ck0aI7Nh8EqNMVv8WZdfIycNQiD4ECGNcQMznZTO2yz05BnKEtyxquUYmcYgSXaQCtRdCdhnMB
q9C2txHnWsZiM7KabEKjp8Nes56bwjSSEdP0zfEo0y3CrH/WW2y7AAFki+U7Msdp/eCjBYqBWzck
18Say326tAXCiS3eF6zURaoHnzw/BtAWYnwVNuAt4FWJFf6qf49TUq3q4MAkxRA3N4LBcvOgCVZY
mYU7qpJ1ur4AHNRYa0v+pDfpffVhWtC0/MBVavP+qrNKKbCgpgnGnMoFcK5RYWPD5V4HFeRkIqBP
ZKvWjNlQEMXuXT0j2I/WGTuhGI/HRwyj/xN1v/zt5hhJYJOGKeDwjGPdNVxjBMqtV3y93GGqEkp6
TmMvrKmNaUardRzgzP9gz5EuUjOobCxnxBxwdtFky9X7Jqld8SHE1C7Y2XaCHdzowBixMRT2++2I
M5vumRpDo4+gYTUyNwyxBJfwQabd6FIXcfecDd00OQ2GoVcPKYofDbMZNQmpmPplMmWMl3HYUrLp
5/eiiPA80fBwm35WL5N26gLdfDtP18pKimv/l+HtGZSFQgiVrpAHpFSJE2nnOYH7I5lQYkGBXqGi
M8nGQpKDYFRyj0NW5zVyCbYuFmvLNjipU4hkTFLfEB39NbfkmFiWjVRCU9zXxH/UvE9RyWMEqncq
MG2aj1ocgxcUAw2Yz8frfj43Ps2mzqcyhmrKWAngJVTN36orrUusPut7MOlzJFMQhrVPkVpg+Ytc
Hq9wGvOnEsqF78thz1zBckMab2FW+DNiOBh3kO7WFvuP+ujEStVz/ZLNJmwsJpcnboMx3HHQAhF+
jzD9U0PhHKrvbyDH8h0WjbhI8JVzDk5w7QzdB3/XFyeD3NaQv33o72h+PQH0ZlXxjAlY05Y/XNj8
WSwmHFO2+BNI7lxEKFQ+oyc3f//yIXezDUnnK5skHj4bXCy9TLppjbZyX77HYrbONxFKK5uFXlN3
Tojh5Lwq+YbB+Ij8DDa+GQMO4CiJBQiBXhy4wxvcCtk1Vs1VcXINABC97Q914PLY3SIeKAMct5kI
igFHC+z3njUKT269JTAgEykXVst+e+H1yeRfV+y41AINoX39YsVK15Mv94ULRcdqOLlR9RkGtuTr
M/kGtNTU7L11fPDFi7sUXE9W1lF0K5imbCd4aB9mDlhGZGGAmwYzexP1ybnaH9KcazvtYXjbBqYS
jIbs0Xg0wIl5hFRewUpryXABAuosUAaAr6sZMxm4R/u7b9G/liXNKWVkWGartklU74PJS2xUowiN
Ah9jNk4GNsGvleNe3VuO7h6Xyzx1APCSqc5FKqLTWkKsXvg80E9bsfLeE/Wke4NF6nisc8FJHnfY
o8Ehp0oSMWu8TwAYmaUHqWN2lmAHVzbe/3tCaLsH1+NJe6h7qS7XnAgHaG3MPMgSHYPRaTSM/c1x
bunikK6sxTBqMrhhDYmcb0uYX6QfXZBcF+Bzof/xCI+EtgZPhP5QA9MRDh/gYfn2QpPQE29Ig5M1
BtQLxg7vQRFpdAELW3z4UV50bco2aXMfdZeud008VXY1o/beRnFjULhQB5cxxMXoyJsUtMee9pKK
TsYZlHyBCbwYg8mm8ecYs3ARP2llE3i0XLpTs1cK4QhTFzA+l+44mfwDxHw5t5sAg/vogZAxLGJG
oqxGX8yQJLuYuR/W6Qzgkb6x0ZnUBKxINHU90nHbJ0rgRSuNd+2S4qNv8pEj10PR8XyO6/bUiJ+c
fhY3uHn0oUT+B/YBjn32z42w2ulfS4ZRskwAr9hPfGq3qo+FdionrbQTDNZ6IRMDBSF9cBwn0a8m
+57Lac1pSmo4ZSvQ9XdObCTOgsGnd3j21QacFhwELyZJ5l256UpsAvHg+FnTzP7LM0DGmlDy7QrH
0kybOZOuC5lPdcNebKtAbHqAbB/ijnFrXmvoZdGa6cYYIrehM7Dl1Y6cBRVmntCUjByOtNNqMZjt
vg2ZO4Onj4OdvhnTis73Rkjk5kA/bLMV+CkABImMY7DZWdS9rUFiEjrSsHUThT063Zop3bEpJmX6
qan2xg9QEDZ83aqI5jZ7AjmHBVCjtqwBgvsqUD5tvbAoKqPJwYfduzfGcXym74JZbmLLDGYO77u2
xNb2HYM1CJ585jbOfejeeRIgsqP6/QefyR+5mQ5ILvsBtbQbZwbzHqJ1pBtcmcQ4CRASNDRFyZ6J
l6LSG6MBgjTqOqyCRv0XRHME9HYqw+uo529wTcCVj7bewgUfEaQMpThECYgv+yZbEc+7NE15ZHwX
g8iI0UEsgMDvNzNGjrQazt7rNmkXV7/iDS+B8BTCdWgbjFChGiKMkpc1L2mI+GPq+k9jEloRRxsa
wNxv6ov8WBHcVR3MteobFQRWG06Q09nTrO5ejgjEq5hgpcWr1ojcCbLM/+vuOQlA7QQXcC6Et54m
GWJov3SXtR7r1iLLC9nI4czVWUOpaasQQOsqnEaXErq8Dh0/eop/UAbeToxzoMD579My2rz2DNoi
P4MbmSRFu+2oERueYokRty02PnrfmT5JB5Ru5m6DeznVrsOQg3umLmp51C/RTP3bldf1OvdAxajq
B8+9jymoKcx5gGeztQC/hzIhhwOUeouYglhogmHkmuWsu+rVLviBA61B5HumTjvWQTxmcZW1hSvX
uRfQYb8RkNTkEL6KGA8shOWXWqFjjpzTgCMcoi2oDDG88ks3kKWtZSUW1dACGBIdSZIzfjG0Jtc2
nxSATYXK7r3GcDCJ9t54X+wLZQ9YNdqQ/czCOTKN+BqHZXhDonxlMDhWL42dmKdQlL/xoUD58LK5
+SbeMpN0bW87KeFlOs6bywBx0LQ5PFib6AN9X++5ejTCF4FBnWj1X2ynTgt7JKVyqp7F1ZBqiB+l
psnLH9+QxJw+HDgdqp7RMEdwwenaui+CbPdCt+Onq9RQZFn6JCaO/mFlZLh5O50Gkvwo/ldUJkeF
EYCEe3VrY5+X/QqJ9UUAqeq/9Lom0b7DtNKqFXkSk4dYEy1wjSXw8ILxCay7K7QmuH4GkuCP7f0/
5j4WgFg0yxFotl7ihnSAN7+SGu4gSpZZxUgvqgtE7bMJyZWkwRdaKsJa8yrny39mt40qkRIheiyy
avgraimURelVQS2pgNtF1AXb8Z6QTQ0BJQ0TVX3RuYCW8MZ1hkrZv2q+4cG15lpnl4maVWbzcczq
7zVz2P/TvKDB91EO6b7dxGs3JdFPfjs+74x4WKw3WlGhF0y3b2AIhuf+nFgkI/ipvCNZH5s8LCzQ
3sdmIM44OzWACCTvtcw+zGzz4qOvy7r0Ek5yAOVrSdho39U2FawraInylRQuBMkQriA3axtvCtrp
FhUwNNzI2/R6fS6hjcYw1n+iUYEjR4+qxCJfTFS/oiUU09X8q5ibw52955pUeWsMkqkjHO/UuUfg
AoaFjyLGeSviJ3vNFJvcYW5/2MaMjTjBl1yx740T0jiqWJZlQTOq3Eo/mHC9r0XFjlZefdZtq5wu
XOuA18BpXWpV6x+hTSvzI+I63j3JC2Qzw8tShNaV2RQmS1hK/B7o+v3PhflBjzQPieqD7x7njwgB
nVaEI/v0/ySIehNcOAME8WPLEGm7jKhd6hFWgvb8GjPG5TCQUoV4RV63Qc3yDduCR30ZIQjiQmC6
dVqAYb5z9ex3ibZ7hJ9+/wU10oqnzaChlSNJpW7s3bNNem3NDE5qxlkrSAV4xHuxxsrpdoJbL9S4
OAKgq6NcUctYJoalP6SzY7dDv0mO0TomzTlMdyIiHyQoDKDr3zhoownNkFyXnO3hNQdQxm+sh7au
Wu/gY6zxQpat4JhBTuNham/z2tjA9b5eAtoOw+Dqj8NZSqkWeIqPAhhSJRiXnCcHD4u2+GraP/DJ
NceUMrXnXlo4m4qUkroCrr1+1lTIgsiHtau3MQD2cIy4LdS+vIT6qHvwQdBV4Dpu7goLwuiIsXSg
26IRetlG7/OcTd1U+3Ccs0pf4gaV1C2Av5ZT7CETbxvrQS8Inmqpvot6JNx39UEQGgqDY5zgT0Be
dvc33s+g9TlB7Yp9f1riYzX7bIJMgUuzitBGzYaTbyyO7jVp3BCneiTHDQ1jziwT9KuxSD/Un3a5
QFctq6u9IfaBs9JFEQenwq3ixliANeb+zSPmz2qb/uUUoo3d4gl/9fUlHF4qJRnwDSBk1tcUfxzb
GsD3JJLPZahuniAZlCVpRHRwkvAEm6zi+6OykzT5K8K4qNi0+qnIPWxbnbddP6SfvPyJkTOjULDx
M3y/wflZQAr3sSHcg7paaqVsLm/l2b2mupwabAOV2T+5aA+H68X/Ck4v8++EdLlQC89MN+QaQnJ+
eMV7qfGXUlWXR+GZaoduy/wC9fN8rj5IHlYO4JoiZY5pwPyx2gHPl6QvxI+EqmnIfg72S560P36O
B7TO2JNVoxuUsCES+s8xx9/wKENZnM7jwrK/Uk+S1cAjSC/FpZqeIAY4Vajd1N9DNISNFVYrczpZ
E0PNJs83WJEgX+pRZLmst+vMeJ1wdpV4Sb+KcoN05sCvl1XPRDUG1wKb9HU+iAMplIYulx0WO7HR
KUmjb50HKENPskt0uiKuzmHVz4j6MGcL1HQsiq+Ok6amSVFgjYsyv67rMxinMSdaBTre3vE8RZxy
JI1rYfIyNfI2VFeRDhGjr5xK1wRpwjLUxEtgFRnUFXTnyvF9IcFiAyldlkRrkBA0/ewNsaLkVt5x
urinrBihGSqqzi2cqLJIgsJjVSEIWhSzv6uBZZo5qN58DFK5IwLrKpu1jqD1V7xgRlrJXD7+PGHY
rRxMZoLz/fnsVVHWWcpc1ddwQ5GMCYUerMW3/HNirIWkuHL2QmqCQ3sY6VyLpN1K72DmVcuX0/dH
lXAHhe05Q+oJgt6BgIM7s1ipBX7SKcyMq6H9HUMK1J0+i4SpwoQsFNQ2ibkhUCnDc8y4n/SxeRGa
PMoLsWlTQyh2VBlapexzTDoPSBvdCF0no2JuGxgEBUbMkl45p7NMUh+2tFjU7QErXYzcv23j2Lw7
1Na0dVpl2NseMi3R1brtyFTfBaIaeEihtM0G0w9+PNS1d6lFjJuzmWHdWXsFxvl9EgsFFjiaVoig
S2eW5coVu372hQIexCghDbGlukbpz1YZVxYWFV7QTfcLVrQ8l8YsxhCtnxdvxmh8vhLRjd7mzSKK
3+USm5Zfr6r8Twjb8R2tJTOl10KKRa8K31dhE26iPNSp8cZl/v8F0MPX1DioL40gXkJ5OrEkNU6w
NsOg/8zfYwQysZovz1zrNFRq9zv2ROTUcOJijhA005+srkWHFyuWO2Ce5eWicEp8VCTp0PlwJTbB
1n01ybw8F4PTNBjGvK7qXibatMjiGtvKAuOKjvb+rWX8gSjRDlLPT/4Kno6RBs104uokRWg1Ri+O
ey36m7i8PSwDfwpbvmfi1wYRdrerrdIFmgE8bEUXy1j5okbLYtqvDiftoEykRc2uQ69rZZxBBPJI
rcXgXJHWVKFJZgcJCOm+kpAwceujdEwTv6kr7uyAAFyzw96tNtAiPJ6Ix7Hn4WRmknHe769LDANY
5ZQEKlvklyX6ndvWjNyq/Ycsl8pcIPX7LqzHIlSS+cy5eorqpjuH7sj4W3ITiR6/kJdUkErQASNE
cQ/y6JmCI7Oz5uMF/a22qZd9U+0/5uKQztNfd9ULSD6xSQ9orC1lPr7Y3vVwNVhAMk8lL57BCgE6
JJMOoB/DNiA+IiyjvJHEE7VMbpVG8gbZM4drz9ob8coxWtkyyXBCV8iQP9RCb+syddAo3M1WMA6T
q2Fi1RXI6NmQny0VsIWr2YLcIZzIrPv20sbPCNyRys1p8YIbLjUf25PlsDtjyR5YZQ40JlLnpv4h
uMUtayeoUQURc9hZ3ngCzVmm7M9HWiqJ6zYkz1RGIk4VrRy2JwDUdIKvUFFyzuBn1ozk6ZSnEZAD
OGsAsOtHRKhdpClLHn9PkDe3I8sFHZI/sa4vo7r3W8kYFXolaet4uMajQzP8RmsW1ryNFgjtg1GD
9bK5yb7vqcJgIpPR13KCOA/GyrWH7N51QIn7RMgaSvGMvSwNRiH4XHLYlP8PTIj4OQHGx1ONHX30
uLnIUZFBirBi0ypOxR4Ap1ma/5SZYcvZqci6d0QgRd3NiNZ6/W9nI4zCa2y7JDW48UtzVGWKe9xM
4B73YxFw/3UidldP6BGTnbxynDa14HXCijceq1qkJ3ECwFT0g69hbDguF9C0CtDb88ntxELB1RXg
92F99oiQsdTAdB+wMWmpRtqezXCClSkj5xbplX6xE+7KNkjDJKMyBzk51xzdymGPBS51zuwktv2k
2aWEHYD2NCgrYBL4mBWE90d2ZnyV+0ThRsNiSZwnkrSQMAExTKmtbR8K+hedbqXG1lFJAqjm+xH+
j6bHDeUN0mCt1aFB4k+zc00CZFujkfYmUcczPnNKEi0YB89tqiTCKvHb21OIzW6vLM13LD7BYqFN
BYeALi/4mbmUludi5MgKPIvjK+D0SDtoMuoad2KOfA2CPLsgO9LkpY/TYAeVenFWU5T8HF4CQdWD
2xmY/RI3WBpO/qascrJdC/7AF3VdYpucN+/qp5IxoyPJRLQkXIEWhUsjGRbteCCI9l6jviOBe6TV
iHejtIeR7K1eY2SBw13Aj4w97DEutrABz1AznGJxgYG2PRcCFt27RuVTt4ys6yMSip2gyt4TtwZM
GvQNMQJJJtdiUryKaYLLPt1p28HI7v64gQETwBFoXFTbTApc7DQoaA8WEMY87aV04gxiXsxk5iQ2
q8NQPllSl5qWg1pqYmjuHDFw/io6G7Zctl/GqQks0WlmaP/f2vp5nsy2yWruJJFx0Jtb3+DPWMjQ
4bi9riv9BXwmZIs3g43ezGWQDbYDa88sEy87TqRZUBWXRznYa9m0n80l38Tb58mCG9MDQifD8i9e
YsPbSB2NUcybyy5pfuJ8wjhjeQ/HiQEhjNH4bYAJ8Nq2rjm7bJ7yuU21ZXb/rOrg5QEi6cDoy6dL
My69KmMDaZ0D3lhV4MWq03ktT3WqPXwaphJYHM2ILL3fC+tgqHJJa+3zyyLQqXlB56ry+IypZtFx
Ut2t3zSTOZ6TNrmlTUTNvGWPELq2+sACn65BilYSDCNtQbN8A020ZwUTUHoN583MuqkrzqW1YJNq
+v13fNy+XB1yIDalkroW3BQKlzxSZdCCGPtYO0/2bpUlvGYGM55Yes1AYJhqnb9YsFHP3/HtH+m9
qF9P5exuO+YjQ9n60rK2ONJzqBI1B09LPFZKI42eQig+y7fz0sGprXZdmBDRcUrLra2ZEKVsUiAe
ujUjF0NbdRZCbgrxK4rYlaSZZb+xM7h6cNJ13XCIgvXUyT/6pA6GFG9apik5llAkrIF7GjYBo6qC
6wY1Qoo70tEGqkczPUvTfMgFHFtQSCTAHmtqQIhetJYCnT25ivuU7EFOBpVOmpaOmWmEFZvwhdz3
jMndZxBpAEL+HG3d7hr0g+HpHcGbAzkUutVG49BXmbUqSc+byPp/j4FXj5E6KAmBxkszA3ApwjqG
PXysVQbMy/4mJnpxJyiWr1tfcKlTvG4Bfv9mcVkoxvd2ok3Hr4m0t4m3jAg0m+2Gsq7dWi9DXec6
zY6vaz2bNS24xGTa25T+ugR7RhLTAs5ZiRKF9SfzM6E7Shflhe6dBab/wvhqry7YKDKJdlrO4pFA
R3ux1xO0iw/6iBtQRxoXYOm0gKTiOL/rbdjV9cLnAJslzC5hDXINDJGN0a+0dxvMioJjHFR4/PxQ
ZSchAanoSv52qareBTxLdRkYkyeoH7jMPIYLFBgcy/aR0Kn+vY8jt86ZI4JmDZqrNfTsykn2poeG
BgvThl2vL5Xp2wOV8A0UhCj7xf+Q/ZpRZbpy6sinc9Id4PqqqYq76xlu2BfUkehOY9CV7smajvlf
DmaMPBlBnLwDmK1AXagUlNqitxlS2l/d8iInGQ0vqndmgYBboAJaPZ3vr+AI6vpVZ66Q1PIwg9BF
Rqc+VDWgbA65UIEzbjvafs2K1+utZtFxhgIyTuYqr/wupAgLDYpt7qLWStflwmlgg4FoZlLT9Mij
Hm/VO8tHi+/3YNPfgi4jAEA5K+PdVww1uBLwSQQ2iAnMbvyKObABR/qAEuHMipk5SLxWFyAy/aRb
cedArooOu21tp3/lcGi8PJMskcsOdl4onZSp5WCcObOu2iFWhQkR6aZw3HXcgrLXLERC+aXQWpwt
f7H664GqJAM5QUVJ6I1JxY+6v9i6xXX/JgwLdC6UFz7+BISA86V0y7rtG9CBuwp34dccsjW4rHJf
g/gpmrRumEpmmweemen1YcX/vPDOohrF8NJVQfPIdPw6Dzo4G2j7SVDTwiQenObclsTRfnZHmvut
/qdXdCH9VNPiTJNcmQVkwj6qo6uWwNsMm/oX25CgaEpLp47kTM2kq80AQspvZ5Vo5wfuTZJNzU5c
DoJEMG0A0CLef6NmfdW1r6eYfvMWioyQH7Zd/tfv7KB977a08Yqi2cRf5e5KD6PJ84Z8gwt+aWkt
qoWCtkd2uM923+HhdPOrpA5oD8vQvE1wAG7RSUjhqnPM2vsI5GkQM3j55iL/bre0i71g1aXoLQfY
bVg2/mlzCTX9zpw9qSApWU7NDPghjNImrKEqA7/yzNKd3hRLMCde7NfndNOVnCtbl+AncsxxJJAm
YVOUm17+i5ySVSWmzhk7hNIL10zbXAJ+z46oBGvJ1Vn/4R6NjXpJnBjVCoREQk2HNTd+0C3k31Rw
8TcEillk4/DVXohsdaIMkjWHDPqc8kGsfmIRGEBoC5YZz0zymqH+OzBrHyYya9VJSALNo9YsWnYk
dbEj05ZvRlZdeelXFuLWedoTdwYxZkza8RzEA5j4zNDIx/mJdN8UFKsM1Ksdi2PazF6YrEg6Dqg9
Ydq7iUj7AeuTWNPN/lSnJ4nqUSANsnjgOJ/rDRVSg9Hx2ZV88wOm+Xpp/5Ka2swk7KeMrfAoLNLb
qUzHLEM4gT6m0maI9gn5CHuJWycS/HOTX8HAxprtApuJL00Lr9S6MhxsITc/jyRxG9OAJOtPkLIz
IcVJMRa8RM/3e8QmqvgBVE0qBNv5Smtd4X5XiLKb75p15WfIFf6tKnJ2y4qbYVlMz54dq03uAjvM
TE9D6xoFzBfCdSUh06/p91x+WD70OBl/+g3+uI0fH3MTrVBKiL9bz9Ub4V5fNRFzJ6DY9HIK2cSO
X10QdsD3Nbv8qNG+IZHe2ls5DEc/d3QQwmegUN8riHgr1WgJMASExzvrW2AARX3ZRgdiudKFwZNQ
PpuNGJ2wpUtbVFmcYejLzqmKhG7zJmeVPL/wMCMwGpOZFOXDAFkYbSK01sGbC1VUpbLWxton65SX
iDwEsIJDjZPunWxvDJ+tJOYNgmL+ezWqz17DSHDYw5bWcrNlQ0XstDZkUUx1q+QW1n14F7nP2YzH
ZfproKNXhr77TlXeRhril+9Tvhx5DhC/4umNJD1h6xAMYL11wPLQpZmXtL+S/QbFsTPr+M64HrKl
5bqTSpiU3qYA+T5/sInRCi2KWylLW++8GO+CA/AsgBSmAE45xEoOj+Fu9ZkVEtgkl9SJYXwVEFIb
ZoMcmV0v5lvi4bxSx6ljQyN7e0y2ePsfIYt/upO+MzPVQ2HoO2VaN2hl45yHhCJE5OSyRfesIbGk
e/UlgWEocCXM4xT5FdopbhNJrp7BJydhpbp9XNibZzZREIbHuQw797X1mQZbsYkwcRliXHSbZRP8
RYOubY4Ko7cjttRImDc8/XCwStz3eH5HC+ALI8qspzIutiFNZ5vPdLIXpdpvXwKnCfmTNKYrrVFv
BKrpZ4raIY3rNGs+GFz9xrQCdCcpmwh6iI3tQE3CfVKhKlpBzj+mvDvfYr9b303BCliUAw8mOd4+
J8oFXCqdg1VJbOlE0FJAjUDZ0ei+fUGaUez8VmgarOjIkAoobEYFERu3x53oFE+/hkaRKteXcn4V
3+eVKCa2CaBD0J/8swYfPTKTmTP0mXsiXkalVb4N1ohqx8oJJPSRIZqljFoGBeR6pxHZyD7Uor5/
l0y4jNgyi6gepnej09ZS+MEHSPe9+vfUsict1AM6I8Rilk8aTHz1YCgC2T0YX2boLW24A+/5YOtP
rRcNRuY+tMio5jKk0110iBZyTajMeGdeJTE/W5Gcs/FqjzO+aBedUzDcaTiRP4MgbKlZZ52DKJ0i
Qcu0BcEA4O53KmefyjRn0n1YdrK8dqO5zcK2eYJr58zlFr+3kJ0WyxEM8FJQwjQJifNpkOujaIaq
j6pTIj1m43B3H9Slvpr+RRpmt5+7LX05piBI5epLmgR/RczvmC+PYGeLmI9/X8DrOWULJR++Yb5o
X/UL14lozJBgvxIyXmuy7Vq+KbkOqCKJcNkWNPOeas5uQMm8oskRInAGGZM9bwsEn0mERQ1qYZwd
sdJHQM8hKv13ytaYQ1gfHxOTo3h5Q9ROpF12wf+tWYqgJfrYfh9RV0jpij34RU2sYJNaC57YvyOZ
Doxy6aRsbp0m4aEadIesQangL/4TdTkrgYikqz3VlmqaGZ72E2tIEaOZaHpzCpJhTFpeVW2vOL3w
ZbiLZOPC9GVLtl/EltEpnJf5FVssqqW6UnHDO1zVIO3Rd/zeoQzCJ1hqU1g6M9J+5N7dcj3E4pNZ
z7Bit9Bo3YmH0264DFuB7nmEY5ZKlEgB1RazxJqxTwhLR+JdSYip2ib51Hp/6+KiJasuupJNhwZf
eV+j6KeeZ20k6mSQGLYwFXo4icDAP0639Hn8KLLi50qlSY+iSU9uPLfHvldmrokCrAo9LBBWSjZD
OUovd+erYsrovk4odXhyZO5Ze/m9vBGOc0avM3/vEE7LglMExVXEisSMsaicbYXz+dng3A94MX58
d3cZf0MTvYm2O2zvD+bhrdBhDzXY4RN4l5MFo8e2UyMQdANdtmSoD1aDqOdSuxOpZDUvrkBzGfor
S4IpIhwPmQh71YRveN9sa3t3T8CmLDI66GsXvKfNcOyK3+UBGCuWWrJ4WpHzoXP1g81MyHB/NVvy
EtqCqmCK/sg0i+C1i/vv+7N2aAfduC7q/u/AIm6lJNN5/HjWyIhE7hHGiMjh2JnXjEC3rGjL+wlb
wsLi0AUdQ0mMFmFGGV3xU+BeDR6qpOFL8HXFEWzvgEvENZ1Lh3HkCLwuLaKoPn8aoS+oigOBXMsD
4fRBmkKIMYkxbaunraYgQFA9fmWeK0uy+0Ww294ruhSJL6+GE/I4/GyE0Se+ctzww9hFudj1I+NZ
aN3sCEn2cBXC73vstH5iXYjCYTysbgj77fuxmKEM65A8xuj6xbc0KjZUrORRHM098qBRJiXAIjZi
aZnwFhF1EvJRLLQIVxy0Zloo6SUIpc807p7zfI7sA8vLjtCHF9Uj/uqwG2R3A6fZE+vbv1+ip8WW
sxtMHmGQGq0GzvnLnopO96nG51YEyYgJ1fK4nxVFoiC5I6P7oqEr8AwTEhSfUMm5iCTAG3ZWKfPX
VZRfGr/hvVAZj48sWNcr4WXYPU1PfZuUq2GobH8p0u9RQfGFXO84/iEA+7a0xA2Hy2Bu9O+0sYzm
bBX3mnd39c1gqPAtIndLjfRrnkjuXTxVw6jEW4hMum0SE5YtyH0BdJQAOoqxyw2fZ/PZrr5bddxj
ZcmPRGg216OuW0SfeqfHzoKXFd5BAQmxIF4Fwcttbco0/xjeejnOsnIa0oEf5SqvEC0+DzVkTDZz
A1uH/XZhbIRt5veIUMiAS3aQh3QAwnG7leMyI5WqJLXZIrDxK1gwuVR5q6HdcC+dPsvSrXbR/R/p
uHSQQmKg6ZAhmYTvoXA8hzsJ/l1bn1YQIv07vG2er+OdJ7w2MoWhhzEKhl5J8TI9Cr929KqgbGFX
OSclOpeYXRJ3NN+eDrcZjoueo/WbDATWEZcMTaYRsJp0tUfgkjiXNlDyaYQ1DROf37p5EZEDAIO8
HEn3OLjLtDTmXt2qqO4zGIIA8jO8NKsdmdMZRPDbSITBsWid1z+VEyqDHA1mfltO4CCLDVRuJaHS
7odFNbweSaTfTdn6xWQ2DGWTMtxAKeoMOgWks4LlmKr2nMUawg/Z3qa6bcBlGCtAfLitE068clzA
b0WdY6WAyrAQ4nG1pIMeBxQg48UTfLPbgc85AFTmujHGl54RlFDlhViMaJhtcsOJd2eRxTDmv8Cl
kyJcxKKiY8DRjolL58LG35JUm+WDPyFX50QEfu2U0QFtyWaYqU6wiglUCtdKxpDqS3JzSNkqd9Dk
5QTlLNsXhEOzfPOcIKL+MwX3B534lK8GWYPpQHnWU8NMcQQNiUw51o2Sl+9HLKeACokuHhjEYOIN
qmScbnnqCMdwA0EmhcVoycAGqTJRAOacvqdTowPJzIKgrBaMGZeFk/2d+fdjw1N8XJoSWCaUA6ru
3+tXKLf62U/g182o9tnKyoGxvJJ4Rrb7FFeJHDueOpR7T14iS1xVE4h3gQdz3+MJWVj++4s5UOSo
Nqj7uPjDbMyQIArCxZpU6OsB6z7t4QpiZXnawwUj0oWxAv+PUvzls0Td8MmYjGc8jXAicHxGJn63
4FGqyd1npFsX201jI3+7RoETGnikc0TSCVGL+KWHKu+1YoDpT0OU7ICw1wpQKaiyxYChHr+9XHcD
OZsSfVA/z7JStTJaU5pzjF8/K+nHudTp8PvJzmRqwkzM60XUsvMAZ7Y/DQ5rW2mMmYAlRdvetASb
xuQSe8mAdlzYi9F3EmSFrDhPe1nRwX1ew9SYeuRMB7Vs3i3qjEfspPY/EDVVJ8rOwXaqxgDbsBKN
81H3PXagHgChaGgWtJMAj4PC3T9Oi6JLoF7fdJh3yGgCn0HhsWMCUAYM5jSqxKtYvr8dqZY6pNH0
iXTIG8r/g660P9jQC3mFzHu7vHucvEjlRLoUpc38vZR1DzQVH0anfOAdy9kr8YraFuq3FNtigVOu
UD1xs6sDWlQwdKfpGPcWOrGdme6G7diqqaWLJ9prwue5bVvaAxzpXLVrfBlNN53rRKsK8jzu2Kmv
c5OUvanj6cDC1P7SQ3JfeG+myDXhz3ovzw5bD3YxQ1jKtHqsRqklywSN4F957Roxtl5ETNoQw3je
nJTsEj/ZrYY0FSKe7cIhG9f56VCzeXu7iF10Ugpi9V/4IbQBavcQ0l/kp5XUUPXCAEV2cMX/wqde
mO13rBZ5lHPYdxmB5KwrBVi6a3kPm8FfLBwbD2p3TJuDdZYlb7eKoK61MSQMMoF3ytD8fgOrFP2I
sZKzGFXuBEeF5gjtZahmuR6mVO/ow6yagTkA/QXutMkPOi8DjIA0hMSdXJ8kO0x21+lpRSGCZX7l
1cNS4iR+uhX6g66UkfUj6LTIcMMZ7Q1G00goFkHf/x6/hOAHyL+G5EpH8mSEYqiaru4ZeA87IjWs
PdqinXNk4yKg9sOvoI6dAjUoFrWPyA1PmsmYdWCoGZwHXYxqPFkU6XeFur7ODAJqk0DKxajMaJga
4tWLaavdbMQIUNSchriR0FXXFlQ/TeseeWUfjeeryrivHJp1bbETzEiChPzWURydFOZOVQ5ZaNed
qN4X3U/0UTax2QQeJBnBF+sWLrIrPgy+kkfCuBHakcq1Mrur08Kme3+HvlpnUaQMJvg1Ol6ybzTE
Mh0bP520WXRj+DOaujrna+0MQwdiHlKLnwSbpR6m1QVMIxVDJbf/yTwfyW21ccNc5s+wT1OYM8WB
SkE/bZ5hZ+QetRUuyRn2OL5oSyErbigW3oLsaqOH9RS/QqDAaISKiC3ti4BFFlr262rhLb0VAEWe
fFxzdXPl7J0dZny79UtcVIM6xdWGzD3ZF7iWn9i0Nq1X0s4dndCS7Wwfd1NLlTNZ1IWAywmQYcsE
NlAh2DguoPko4ZcGdSvwahPMFW9kgVNE8mYtT1KpR6/KVrfR8C4kKT/M0tmPkG/IErLUc0g2wO4O
5nUYi8ACFCXm1DnH/mlLqGxGKdU0AT+W9jOM+Hby16YpDxt8A/eH3adYgbV4edZ9S6mheSjR6OLz
drHXTpNONmOeUeeAAcQV6pTrzzPwpzjXJEY/uUx8nYsoxcnKZ4bj/T+IDh+SXfynXgQEEIKCyyvy
SD/7bcbrZlnF2SMkU5y5MqMtyB22HUvFs7Q+9YYYtBFGtDqZlxzBRMcp2HJ1cqlpNL9bG3Z1aPaE
Qv8bNFJOFeG56bbl1BLTF1afYQzQJUFG4YUeqJ3ZZBCBRa+TrZjAPhhfBRkqMymBxSYE1g40mAXB
bQANGCi+Yr5YF97PuO37C2MTVcHIn0SILWA24ddA+B+QRR4HxRqfQ31taRnK7UdLLfMhsbxxorjb
AGghuDwt4wK9rE6My3q0d7ei3kYB6EjlA/Pajv8MDUB1s+6AvBHI3GXNOzZWNN9AxkodUrZ3w++B
o7XIo26zuRTq0AbGBjpcczlRH+3Th+OF12rO9CycYpf8JqsyhBL5sgPgRQmJ8xxgazDG4XmYSa5P
JDvHeGiy4MbGrL5s3v1E1CNw47+SehMzOT+aV0x8lsb8iNS9GKjQEXeV1huo8KfOlg5Clw+mwoTX
RsmFY41arree2MxMN2lMWdEinEzmFvQi/Xjy9rSa0HgwuX09hwAloTORhspxSXs2fzJqPRnQdVUU
0X0EV98gy5sV/j81cOAgxxIiuGjLpmz7x0nGQpNAQD3blGrI1vpVfeD9xYAiHaX6h48FTgSWE+7e
1cy5fgZoofh2JWCWwOPI9zDVIgIPFxiBs5M187GADwvOSjORLPUgdOQjbku1zAJ6uEOtb582Mjim
ENKt1gqSleD6/Eb1waAn9uCxSJQnmM3X35YGL0ko3htEH4pLc5gVyAMIKFUbrZ4lxCuQClpsCEzu
v8t8NjA3LvqqXY7hsFZyUPf9hri4r3lOKpS2fYeB9KcZFC65fxDJsotoXpf0cy/KAsqdm8ELTqc8
0VDi4QJfpJzSalCQsskXyEEfSr+Bi2TwKobRgS/jFHNH6MA6lkCsweNvnb1C4x/UXjL3lDHscbBQ
XqlGTqMKbB/QBiLRdkin2/Q6xL29KMViCMDM5IMQ0704SJgHO2k9xocR/3s3kafKpGZBUJXNnUeG
4bfQrDUEW2rvm0BUpHCinxLzzu4a2bTIDYU4LMOrgNO2kujho3FZbVlZJIi4oPoGZd+K4Rn+2Fvc
c4c3yrZJuW3ad4PqyazPnNvBbdl1C/98zYlkHtcYBK/MN0kuMwa0yh0Xz3LOc1kX1eMaIMg4sj0P
J9hJg5+X4LvbPvfp7WIywQ3uBGP9x4FfRTo6cnD3CGRITSgcT3kKk51lgmIMj0aGa7LE0zrQMMVv
gMiiPgvcAQA41jv1xN3gTeGymhjCRs5RTTwqfgpCpC3QMlpDHkjmTd+nxuV8pcJt3a7yQkD75uV9
boDpYPYaJStQOh6VBvC04TWwX0vzKBYma/xk8cCYlHqNtwXlnlYNWtQOB6kE6m9PBAKiJygteYIb
2InnhzudNTJo14hN4LKRkwj03TnIoA932Y8IM4b8j0xgqiyyi4+9A4aSuu4/aJt1lvvsuXZr5qHa
l5f3weVBha+IPYUT0dO769O39eQTHt/qxknCC1TjBVpEnRLahe7KFIgfvv4FKAY1upgcJEPrWnsi
vubU43gaQAspCZblULKxI3s4Noz+4/oK3i0TgM1GNSarl27AyUHH+grbkZvB9022Zw5xfXidRK38
3VOz2rTkNLJxMu1Eanu0QvMtLa7pA3AbSNbVojaqZ679zpUQLtFNsUIcxi6igVBEXwP1tWQNerZm
Yq77wPsdRDVRPxEkIiY/WG8nWoh2xNhUE1ukQPmNs8qzFRaPMl5VMWVjSP8/GZc8YeZP+6ym+qcx
xrI0kCvA3UWw7y2JCwXBAxuCoodLIrgBUCjCbgvp4xEwqX02iwAbHrTsDuiw8nkAZ+5lYBtKI3LA
dUAVEZyEefF8HHEQiNl36hA7378lTTzsy0UR3HqeoINtYnAtPmbRKRf1C3uuQLobbsoN89DvSzpN
7ZBc5IxEYsPZvcQGB0NxAQiiRNRzncCnXlku4pbS8vRFJl3W9raMPaS1iHcJ6ePFHe5GZSSdqNM1
nPPg8Vf0Ortdk7P1Q0MacPZtgEhd7vw/0LIcHYUwQ1XGxTmQ1QklQSlsTokVwS7hiSMB0HTA1Z4h
+h44xllOCj4uOPlCocVTY3BHtiEcFBYaBGvDiDIkHpwPAJaAi728tDhGAQfUvYgECYpb/tKqGRE2
p7DQgoryK2O2/6Lgw05wMrsalsG9xuzOqn+/PvjndX+D9mji1SFZx3717IakOP1FMyMH4sL8zfAH
ZwkYKoZusmmSh/jY7Co1PxtJAJIaJVdbQuwzm3jkmm96+rWYn3Krut8wTV819Wb5TkPLzfQjfYu1
yJYramef7t7hikkughfrR1roiNDxkF0DX63g62Us+9K+ncJgDXRIZQQkRJDQKpgZGHYwygWJ+q9z
9965JmLHz/JwcpJS2MhPLwCYjPoR8ae8u2mf94F0b7P4kApFOyGtqa15D4Yf5c1FU23l/rLIXQCK
gEua2DKpK+3mttaRfhS1pILAWmep+B7eHCmeP2S5/gzCPVB/S6DiEIt/gKHGHdv3sIOirYLdlejD
JMog9GTfp64WVZeEbKO8qnfw0DCTjv1wBJPG4nGhL73pRKkCviRaXW+/tZtm1sPgjp9Oo5BMCbJY
uo9PGT74A3ODhviDffGrh/C+IwRp+iYt4l+stwVFRRdomToeRxOFdGMkRkgSLvzLV2p82YWllNza
5odTsgJHi1nCiw+A5K49niBWvKCO2tApOCCc3vSUoykmRXLfFSsez2fOQbOltKF/az7HRO6poFey
d3vSzhSgR5WsbTkVhxUHhL2EVw/yuRhzbYEB5s2wVk+2jUokcjpkM7K2DvMs9UY+gq5y+0RuhUo6
UVJXhysDecmmvtby5j8G7OD9Ds9X4WxyWHEhWuIZBTcsLgrYH1c7IOf99Cnr8itcLigyKlRyXXoK
66HOmuUgiDPnt48HTxthFBHAs1/z/a+G/PmTuwPR96rvzZ9ZwFbbaJ/i9NHXlCJys48VsGeZiEWI
V+0/R3G+g9yqYBvAtIj8m+NrQMxZsxhKoyYgLF9gVkWiTolVHf1p7Vy/ttE/ADcMBOA3ItpmjvfA
dGeHzD/XSrgqn0XWR0tCob0wRrJhrCEH0UB9+EmVsl4QFeu6q4qN+5gJxRUfATZmaFJW9zFaBAc/
DNEf4dnF+Mfg9sVGzZAkCEM+gP3wPaH27VTnSQx7iHwK3NzOz6d4w5LsbGn1qIszHTWBF4a6I2ex
7dNpqqnJOQzUUbblU9RKGbQRAnAdyy3hoj09wVSK3C0Cx0Zut9dzrlEBnv0HqK2vBydrmkbnk2Ei
PUmW3hrokdOvQzDReazwM5SuSNujfLhMOyvFudKm/vLcVIsxD85VsrcBZtc7C5S/DWGE+9nRqmFf
zYygqfUbaWyV+8Gr4rIMfY8CpEQRoBrIuD0uDPuT5yx/OOIdTHHHlPEEhW78r4FnsvW98kUHxftK
kji3iuuQPzhscVc8q8/4NmDsgRZHqgrsUm4FgGsRxyTQBf7GG20l0GYeNL8fHV66lEwSpznORAbD
FPTYf61Rqxg3mwWIc2RU1ayyNakyFrbUokDZVcvaC6XBIataNtrLC8qh3sN4qbkH3dWBjpSmCmgM
y9uJN1hva3LpVbCgDJbQ+VpFoeqUviTETsvl9+6GvS4oAtu2lhRfyqHhwEdcIpe7k/gl0I+Z1lim
RKjL/y7/7YE6Nz+KUsGKbF8zqr+238EDSPni167IqkqieFe1m8ijwlZYmRMQusLNa/kNUPQudx+Q
v26YjZChptHOsJ9Q6qFJTr9gj2tzRL8+ldxxaTyvp3ERgwWTWpTQ5bMw1c9FzLgLHNewL3e9Z+I5
dR8PQtXlT3fWd3DceGC6aT3dObwPJ/hhZ/CwWG/aIXgNyxBRxfOQRF73KHVTopdOk7gMlDCiwZuP
W6B4UQIFfjuqKL5lfxI5BrJ3MNHnRDeds2VsOXmIcVATz8UDwAWjqzRhGfhlbs88W1YsGzXV2p/R
0uLcpwLz0yo3cHTqoqr2iOB6NCEVm+Q707nBUvSI+sHA3NI121BByphr95TNAu5P59mbkHZq8VNR
7y73L8nN94smpdFDCBWjM9QQ3nr7HhxGk6PUEv02s/UlkvPKJTCfPyOSe1dyvoLvpwNAWOabrY8Y
3aTXzmJ456J7TggKE+UygVEa3jpRP342OSRNjTJ3Y9aFAnHXOGlcQuc+BVBa9hUiKQeOUQVOSYcJ
V1SwAuipQA4/Uj+4VgVHtUTo9KVJMMKYEinmVQYtwXp9MZDDnEBy2Mq0quJDAiSdMOICFtXComTD
Mg+tjhGmxfmit5CLfFAj60AtaQ9y+QAv4ZWgEiT/gijjjMas6k8QxgeU+BeFqv9O3kPSURjIz4xz
dpbqOxaADFWwhfILRxcoI3BeUJjzGaEuOdAzGqO2n/pd/RJrnw+tJDS4upb9xq6ghDYsbZdXRKv/
KnZkCNDfJmj3frWnnJ0ILFhYPN/YtPBpCBHc4QewWBHjkcy1q6ifGsmTddhRLiTg2z4eosCyHDjH
eAjdUklxtPSv7Vg9wEvJxOtuwDgo6JUOnsXgJEWtxlywwCHTl9xyGVYxCaEELdCzN589rYJ19gfs
6z419kJDr6VD4wG2y1iURm+oYkFRbbQ68pAtWb9v0L+DnifVfn59tB0xA3IK6Rt328DiixsVilt7
09xnNhprXrlgswkbDZ6y4ZOrQrvbiUaK7CVRNVeY06XTTbIB2bv2CVRqud9WdVZUpi7gR7HbOXUn
8RIZLnbnTM0XoGuyg/ywvE46YFr9sXeu6sLlM1mBsVzCa+sl4dAMs8L2lJ2//bA7htnZvStT6jre
1ha0s3MmeNU8/TpBXx1kzxUJVYQZTnucdMdMhDVinAjHRdnB3AH+X1fSAt8oPqBU+lXOJeBZxWO+
7/ddTksCtwkDzkkXt6C45wo2xZYkuCNPywsTWYEXwvFYBIur7Sn3Y8MPEvtoEsUL5erEbh5McbvJ
HjPOEJzXAgoq+b34Bdeam6eAGp4zKPZ7+L/6YmlBByTWkYwk5j+ccJC+yRwkQD+ouuEOoeyDCtDO
9+T7N35QfovM+b4lcLUMcxX/SroWDEmmxrA7y/5tWGMKo0z9ILLTbyhJps0Nag6Qq75eiZe5vRgo
gXD8d0bwamSCXuppaRnoepuDFAXyE/ALPCUpVN0/3rhefWKEqtpZ0+XHoY8CkTY+8R3NwVxxwEW8
NSpk8qe3G3RcOhLoIUwTqQFcr+OeOwV5lDchgGrxP+3CgJ9m5tiPUs/a3WDX5r6vJJNh7RDd94VS
7LdJ1j4rxlKIXlrxG9zBn0ERXsVNGyVI1llUuygVyIqZuMmiM3saIaFssXu/ZtdA82yQotS28Y+g
Jct8cAeK2P/cd3aKV89Qzkk0IM9Z48MrDOINWFMQLtteHFxQjRrZzLOhQ8vGvxVaYCatgUGAqyZm
M6dj65HurLzr4yVDQAHJVcRsHHujg3UlI+s7Ylcmty/sltFZ73RGFHmSwzqOA624bNcuUY4tYNch
D9A4YEjp1T6ML+fc5kmr1Y0r0OYWJ0YvoMh/6z2ph8DlSVXzLGqvxapeJhjpFQufkPRSyUT05Fgy
BhAEq21ZFYbcJ1+c3+4zDKA4cGF6iYUiKOhzKNL1WRMV/fQXTHE5YFkRrMOwd0JsoXK+KNtb8lyp
et4X7gaGII9sCiiHRio0fh2ttLCNc/Fig355fMRGTszCb/j/1Rp5OHR8pSa2ZRuoggGBB1d8lfKm
wpjVIjIpoTP2kJRcMSCVfr+ckQ3iEQRuLwmvo3JAzlrmVT5PmteBnNZ8030b4GetQKmTGiDmDNcA
3TIAzEld9ZEL61QxWBJcjvuOn16hcUSh6pQAzjXG0HPYneEXDZ85I2gJDHKmTNTA5nkWc2hCfGUA
2eor9zk+ACU5O+ikU9vpvPgxBHxYaGc2XpDLrADcW7bMkOEvU5s0tbJ55SEFi5NB0rS1LprwvJ1C
US9l6Y9EAAWwoPWxWNMuJow6yKo2N4/Ljl06CtaCG7WbVN/q5Lg4JB4MV0UZfxjToGby051m1buT
Cv07YuewBq1UicRWUJNjCrzBfmOqBX59tCUHtkkghoDXyuaYxj7fdkADRcGdWWHV2THCQSnI7OBK
P2357+PMmf6pZDZSxw8TNUUIdwBpnLlHdB7OiTaWgdishFK8iv/535G/2sAeBgQIZqSMVmI58Ttv
1a16QsZFUkvUE/qDQp70uxhCJ32SdPWQ3t0lKxITByeqEWj6DekdRNuZ8RIB7whF2CO0h3HV9iUi
Yl6pDcU3mReiffnAvJGk54i4RAMH1gYovFyS3NfZiH7zGIU5NouwufPi2hgJDDrT/8SjU/KZsmpg
UmGJMlTH+k14zc2rVjb/GLd/hSaYwgQzNkC+cnEzC8fEk1GLGyYD8CIr0bOYQ7WNsd7QxvdDowg3
sbcXzim5mhayrWN5F6Av54tOu1ZnTm574Ajl1tG5111tiygpTHs3UNC8/JAOZxe+1n6GHbgSVTkZ
WemNxUfwEKRQv2H+ct3OINGd5oxc4fk9pheot+hBH/Q9WATisaWcVmyJwUPJbUEDqNkbZMenUiAa
N2348OmRkgHY91pYAlequEsFgxvIzprhw+fc4W7XdvI9VB6c4fneSQaCZK4/nqbH6ObUu5vvbE3C
c63+sq7geanO3UgCFPJqlz5+nA51IcDYTftjAHXXzDtL38Jo+TDSll577u1gaEJl5RfxzS4bKPpv
HQ6jYjfsfWaosN11kmcordCIkj7kzEl6D3qJAUTjiI+2AHI8Ad6BQMlDSQ0JGVk7for6FbRjPimT
mfcdxN+VrcijtApGufGTm6Is8LtNSHF6+EQ6TeXxv+wo+aEbtHdm79hunBjmCBsMUszkCAH6Jlah
zHsMY6PH7Q9PSAoJ8kFh2HKW51NmGPukZQ4woXjsfVwkHsUKLnlkSiGKp6V9AVA/mQr9l1lvMn+V
BajMkqT7DccstEBJdBqcx26PiM0pZduTwRZY8W0Um7St/LhntugTLreYTyxqdg2ddvzjlQ6IVMGI
YLqqCwanmKoDoGcWIza7abSj+r6Cvh8Qo/jzajxhuNAEqSgZdoyTJWBe5+fIy+tM1Qh4giTv1Bsi
AopCOc8JVpFjAY7/DKW5tQzsExfHWCZp7nrNd/t9SI/0zQopA0Zst4bBrLogG8AIqTO+R1zpZsxx
6PK4KUBg+Xi/VSug7rDZnflmSu7M0k760kb1ZHwRxRxcjwkFLgjdqOvYFk8kF2cuK8o121v8wPOk
//HRZbwJ+MDd2y0NdBEt/0vdGtH5uE7VeVbobvpSRzJ4zXwbs4LPH4heeQD16pwuvhFL5GVPbGWR
6pWBM4V8mY+ud5URMmOafgRZFQWiTL7romA+KAUvj9YuGK2eExhPaXQZdIltQ2IFJfHrvECVcNgv
LP2R09RBB4j1E3qpPdjLIQzvtw2Vmd+IqG6CbPQGyhOoyBSPIGRB5ZYoZE+iqMiffXYtWajF5+Ol
Dqbeu0afmppQViYlStW6u/gvYSZa+VqjMP8JXQrmTALc4UKQVQkNipgWTzukDd4dShRYW+rQR6Dh
82ZUtLudVPMIMtyfFbChcIH8ObQh4c5K/CDapWrn8hXCy/8Jv834hosBQFA+/E9YlrYznJFZ+KFR
tqwAhhLayg+ybmW5pt1vPwcsV8/NEg7TG/+Nce/3eusMmeu79pLsLZySDyf6xzmnPVaTtiJAcBuW
s0eFdEiiIEiFX3+qc5dae5IMoQ2/vTKvUcWULHxJwzegyfn3o7DBJfejZCmaf9kv5deBqXm0xQi9
eY41LohSlnt9uEZHbXV5ZsB3rRAqaOvlNbFKr3DfoBihsz22JgzPGTrhSpM/gvI2zNOEoC9YN5fA
hwMmuCLNFhP4HEdJsiEOZQDzXQO5qEH9F24vLOO+EdFFN0ltHluRRM+z7YFSQQecIzfHXVTYPeCM
m+fK5Q+RXW+FI01BrEm30i5F9gEWVI2HVKMCPl3fiG8zhJpw6jyIFQ2Cr34E8W9rBBY6V6+cdAhG
OETbsmKV50s6Iku/Mb0ZAUcBgkYoXbLQEcNoFeayCzSdgeC2YMdG+uaugEvL2GHIYOmD3C0tQvsa
ARwumO5jp0WXa4c5UuOHtE76IVyTwcOoXaC31cJWS21s/pq8Tf1npPFlnq3pVkxdZCNC2RAcDXnD
Kx16L01wuDfN5bSgukoOxMXRd8lxolpeJbUz+hjoW97qs84WD0Ucpip16R6dy6mDlFNYcLD+oiWq
shLcOVH/aUk+T+Pj+uY7SLQjPrLUr0tOEavknDwjW+M74tw+SdOkew+FzhWZfbZ4upDPrlA2i9er
zfv4Eg+kcFD4ygGq+riIlM7M++Vj7gVk9XHt7Qe2bYtrTIk3pxLOihWrSXR2nJok5m4QOcFTKcHk
Q59nL6Ev4fIwvBmIyoSV8Rb+c6pRr5AhZQlr5dJjHxKuYi65vQdHppBQAHi3AV5Db3tQS34w0JxM
pCwrwHGfV3mAstEB+zVHj5UHL9b2Kkt2n8MRh9zh0TvcoLK9QoF2KRj0xCoIxu7xmhVVbTsdUCRV
h8mdQsx+nZzQsv1s6aL1HWMqlVHMSLu8iupvpk8NglSrdlkk+ZtEy9Wg/3YgqKpDbZybXoDLT255
06vlxYhX7wHfHE+2O2yp8KbQ5hx35Os28SZ2/RDf7JLclOWb35dJ0Vtn8+Jabh/UMZ9sZCUMhTSj
lhIXRwKSbPCLysdI3uGtz2FA99fR61qEd86gR0brPoCB4UbBj/VhPIYmdwK7CJ2dTMyFbJ4dZfqT
vtFerVq3Y3gpAyMRl5wevUFSAACArNFAdc1qaV4c9dSZpeN39NpQVQS3hZrVr++9esHSSiQwWGKh
aG7PB+k5jhj7DJYi/Q7/ff7CZS1H47Zz0r+p76UdVklxGC7ElfxD202WZPY3Hiuof/Jh7UVbGsJd
5RrlZm+VKuwSeXwrs75n///V6LjX5I19xWPOWBuG6FC2whvAIfeSLAptPfa1QxkZFsHa13wKFwE0
vi0jhF59HnIEkKp513W1v7MwZX77yx0qqIzmZl8RovPUcd/PfBXz1rV2gcM6TkmG7dQ4DUCwDzvy
d0YOvpKH2f7IuRgu9emidFE9XeCE+5Yn3p2yS9dmi2F9DIFW9gCKuqnlFCK1i28UY6o0sDVu34e6
3N+D1pMHha85bDZMRCZokcc6s8AMFSvS2seo5WRTK9X52vyH/NDtnV/ZX+zBSqQldqnuTUVHtpWj
mDBedH00P3bM/kOJhymFW5KDfWDp55/5Mjz0AP/ucoaKLaj3Q/9/patSPnzQquQyzq0edVVJkSJY
o1vI3XDXukdlAqe8lkqZEQUojBx49TQIjeONmEiapLiYxq96umFIwMPe0XcBWSOfH8iTI5wHidXA
ZwAGoR7sUOrfPNF6wYy5B1Mxw0M6wkVxOLuPxI5FEX7EYS7slYcmFz+rKaJOI5ib2UE6Bdzyl8ld
vvz732n2oE5dx9T1KY1Dq2eW6jLTp2ShORJJmC5kHnSXm/ydL+qHhdC2b6ceSOqjZf9fmp/04YQj
UrT4dJd+61otMPRoGqbmJfzeGwcRb9hYbnVGWUUteR7tmV56ROq785AKymLU492/OYEtpdSaDlP0
WqKUmJsG3P5RTTpjY/MiWwrKlhvXG9/hd95iWGucEQ4lj75qkzlySZ9FrbTWRxn0NGkLZvhp4GDH
ysL/ATLfUAbkrSdj3p1w3YHEyLIchH3NXRTPbtcotW7ckb2BAX1M01MEVMYStaPYP74MNGR7LheY
K3z+bUYFkOgGYEFwEDwEgB/HlG3WT1SzFEU/DuLD+XDPfdpNQ+fGMaPL7hQt3lJ2/ciZTR2fcXLv
QbItowb7xGMz+ZBxHlAuDS3JMJ7sSFUTsFJiLukg3SYjE48GL+MCbFuQK8cAjd+vcPDrNqB7EyTg
by88F6xx/8wyGZZYW73b/2eRZoai46jaeKw9JqnFhkEzNN+V35ebcuZjlCQn+XYZZBGaUzyQCKMM
kOaXuiDXzdrLsGTAZco8aMqC/7D5OOLc72LzCyZQl4/tby7DND4tIVUOZe0zwKt/CPt8tS9Qo/JV
pyCRj7cUs5e5Dy6AFWRENg4Y00v2U9v0e64knbRSEcPtuRgfO+pktDe+NXiwWGk6G43dvvI+9hPM
qsCthXTCqUWElK0d/o7Mu5g05ObVBzBhp44SaGRH7awuCAPG6V4sGarNjePDAPlKWw46YVivQC9j
/N/prmZkYZRaRtuWqZsOKeq8S4zbWWGpzNuSZBWZEWt48CK0L3HZtj8iCWTiiH74WIMm8OijQ4nE
tTl6VXPwyKlUIKfoLyu6kfgEjUXRmEiDfYaUDTGPigUoj9Q73aW4KasQW76Tnpr5G/PgyJshAGHF
IGnyNIUJcXDOrs57wg9KL5DPEFMlrXRUkqVr9XLeUYC3b8e9H73af3/pauoY8ZSz/m8YvfigxZsr
d8BS6nBz6FxM+iSkXr6bIqTvSqCzhv5kSuHDKv0yhK3F5krCp5nWq9vOuoDR5bW7baCEQRIx5c6w
dQkCeduoRYp7jA5UXKChLgbcPJdIEtF8O2oqI8XfwXk2nMpRAzEO+Wect4gGpENdjLj3V1Fw9X/B
npi4CjfuQHdxXQb2Qc94oUxeV01ENkGJt3Fc+bWmz7vgWJYbGzjYA4cfQLez7IiwYiuM01u+LVku
7fFCo64bOFbSNxeAN8UttdvKgCyroLyZqtDLkPkD3zn0VUwQw61iAaF+imcE9xjFu1yysG3Y4Htd
4MCqx3vkTraCwzBPsbt3mqY47IDhIOAn30LIuQEFHRNjZyqKTBOIZGzVGu06/Fo89VAsBLYGaTG1
KEBaFfNCvvn3DtoSszx8b9zrEEre4Tw/vI5LoilPawLQzpGgnnPfVS5XTgbPjAkSFn1w9rCpqP5f
KZF+WokTBj9xKwpNOMb5NixwRziFucbvgLdpCpfUjXr/AGDjJIse/YiA3kxkB9ctyrsCo/AfZCIB
MXuNunl+eAPUF03Q+C3QRjYnk9YI6pvFerIO2pKIXi2PB/DIzZLPA+yCt9OSynO9UJobh9DZcViS
/MTlX9WVrgs4ek/SZ0cjPx/c4aM9UgAb2YoFfbWKaAmknZfm6E/Hh5iNDnp0Qg+kiJ8uWEWwcCFN
ka/DQVKkq/hdqG4nju5F4/clMibf1T9A6Qh9x/Yn0sh9TeLkNVXm25ygeJR6DHPmG/INuG0XBG/H
Ze298y5yK8puHZzvk+BMMSmUDUy4zyc2K4itH0QtIyvlQrXwfDR+MPTBn30gfKLTQxRDIjVjG3Aj
hh76O9eDWDIS8oup9PkkJyWNSXNYcmojIbGp31QdoWYyBG3QL1IWa3PvMaC3pTdM7nTm74ezuGWm
4/pFpPICvS4RDMeXbrctFeufXzfRQw4KUGSy9Hs9JS+VHeR7YKdw7SUw6QpBzwtsozBdRxndnrFR
AdU930vTdHECbwVrVcdsxyOq2ERF4yEH2IY6tRX7vPrhmmWbymQxykt7Hr/hITC9Ty4xtYYfWbTc
YwEX7Oyw5/q8N5o7zFgIakVDG0Zvl9ED2lDLoHK2aGF31qzyacGd+watMK5eBDCLSOfbggXNlOBc
9hP03j7gqgkFJ8isZuZDEreeNux08UuX7H6WGucDwxx5s9GzJ69cbe/zWrBmmGJKW4QiDJLiCpXm
tzwNOOCquj+O+nyJHO/dhSwYwD4iiflRMYoaP7xGhfo2MR3khoupuyOttxdz+82xeFHwMGUAAlOW
iRs+zKruAVdUuqxlXm2bWDv91wPAgYfu0ckVVRISPHiquNYBX1uJbVqhYeYzg0MUEUyshorhXTDG
2fTt1NWh8/ZBOFaKkoS25S/9zerN6VfLMZs5653uouzj6rSPvFzT/pQTMoTtXxI/kMsQN+Kv9vF9
ZwhKRtX3EynX9qONXsMbAXl/UJFH1vJDzUqgP2Cq26ev63/cS8pAwwnVK1iUcP+sdDwMQn7KMP3D
Y6hpPb2Fs0dsdJw09VOgH7Jea9fFXcb4qdkmCZ4sJXpgJFIHABkXbvdH0CZ55RIyjKGWOO3HFMB4
htgDldEjGYD4jUZbm5uZFjneu6WB99g7OeusKqC2U5ntQN5yLafNMecIadXIUHsFkTbLC6w6LSaN
zHZiy25EQ8B/RBakwkd6cPgf6I7KGbdoa5xyNezK5fgVvvmdwbrrgup1mh6dnnI6ZPVzQdthPXsq
anFIzxyWLlP9HgjQRclYy7PE019+QJvlCvFr1NibIZIN/kgaOKUYmg5jPr8Q4hGCu96rFyf8zOGU
tr1XgutZ4UQpoeznsqYt/kky6i9fBuUizs0NSkH+EFVkWxYNj3+MpmW7bq/vp0H4Qc5Id1httEqt
uH+/Q5HPwWJ04iPZkR5O7zrRP9sfHOJaf44HNFt3ZkYlDNvm/8MILTHcK8hvy0behycKJss+xDtJ
d6n3K02HE6NBz8+SFLm+3AiLNVuFdxvQHI0Oya3owrv15sTakiNPNUbAROWKhe3aABzpdulL8Q1S
7M1ekgsPfqTw7hhOX3lif7dJxz5RXtAqq6GgbmHZU9ntC3D0n6ea91Ks/an8k8qykub7imPGreA1
gHvIp4xO2HCRCWEIY9K191Bj6KEOo+jOW5mwcgHxLgXOuLvLCIwDVpETKf0MNTL4BYFWZAlZnwJO
/DCmo9/2VJyrOfLtoS5HQE2aFfFxVyszExvlFMFKQCmstmn5gzcym17aFxjI86murSLX3P/XwYAF
Sy4HqkziK2Brt+TsDn4V2m0Cam6cBTdXOLGomqApcsMoez5Cr6hnjyVWvAtcxGbwffAjfbIn0Ynp
yMb1P45zg5umP4VmVwIFikYHmmsobJUWKwPp7ysDBQDOojktU/dogzMaLkW4H1fgmb1hJ1aEDopl
NoIX0bBMuDHBhyKu284gIQ9VI3r2qUjKhZb+W+W7LZ2hCY63oHbN851tzWfBHa82D5Mh7GKa9bxz
8coL2AgxwbIfZj4ghbccpsnGy+/lrYfA6Qe0+RRUGwLlyoLWNfljdhjEV4gDaiywRxGcVwVj9gRf
mPqm1zJG3DPAmg19oBxf1szry4x55bExkGc/ZdOwCA0ZAlWvE4IQhyaE47CXimMXhrXOGdjxV4hb
hhI/MQkQBnxP1zw81aVcZl5CG1uw4jPdMzJlD59uCA7L4K+dHOUln0K0VDF2we/wgPSzWR2HYHzK
azd9j215icpozLV9M8Wj3p5YwfSejnddAczcOouGkRhmyk22/qQU804DHrK9YlEwPdnSq8kmUs+U
y5o2nNVZNM97vA1E2DxCzjRXTXH6RyAFXyNPaaxbHs1RCou5Z9v73+VdyJAXU20OVEn5631W6i2k
+Cqhs0nvz9T3Xx2KLnvkRWhOWOt8324bvjXRIzzKu6qGO53Qg6lUMof9X1Umlgjq1Y25dmhO5wGg
KmkDK7WMslz/yANBmGg19AoRhqp+wn9ipgXf0OyKINiwTHGotE40LCQbirqrL6OvnNh2wFrJe5pd
3YrntzN3z8DrNIi+xrBw6SlQvnRW7rG6TSnDY/f0iLbDf0y11T3V4C2ZaHbUijwSRK+ufG5WJukJ
n/Xw8tsAJFgucK+z66Qc+GQrhkHYI0V/9MD1psrJl/MjT7dDRuL7M0pVwMsBsw1e83zABpsJ/pT5
YKWMBmkYQ4y/UalBT3xXE0fcSpK+Q3ef4opecfSyB3MFWjtNZKB73BxnIy6vRsm9HOZGESy8zRE1
PnFiH0FKM4ABzn8pRDw/TgKtvJYkT2ZDaxu/uJc4zXbktv064X4D+GzdqUxZH2ofEp29vLAKu037
/XYfsdP/YdJ92er7HmvmmJt+7MkbT/F7zYc9T3yNnky1aEEezxU5C5ht4CkNcErrHv3kC8WLh7C0
Fmn2lzjvIePUAbB3tM/8bd7xuNlr2qwQZAMm4ANwB64IBdw7h2A0xfxwLPcou/CiUQdYxZBrIqhe
BA2mLX1WQ617gRTd2uXG6GXUXiHwaHKfEWIH4lIrQAirMoeXMFOeuf1zsBqmhMgqsWu6boR/jTkr
ABY3aPJGlc6TGoQGQsXuSpfc9WXavzoQoVrl5AXC+8YC8qmPRE0U/cilrTOjViAP8O2iPsQfmfbJ
d1pQP9aFip3PVx7eGi4klp0ifrbeWW9TbW6GU7E+B+JlBLi85UgJi6i5t7yZ4stBS4zphfSMwxEy
ksczht+2FC+H0StsMtEQaIGfNS4PH9hc7AxPMoECj58EGWO5Bzh20dMsMClJmKevDMu/fiUrEXG4
bzbEIsH1ANn2d7vRjVGGoe0wdNFdOC+twKRVSC9vnV83t+sZojsM/P83YC/3NiT+4/H2Uc2YiQEm
gUIXic4y+VJp09hQjZisjWZ+Vb3LbC2/xyjE39v3RvAjAxFhRFrdE/A5hO8uOFsVKddlsex71V6b
nC5tLFJMU8G70jBHdUQ/6kEuGrJUusdChcPXsRokekJoED+CO0QdQzH3v6EaCJLeBmU6LAAyOgYS
GDJzT1FtnhKLHjYViVcwtvj+aFgjDjUW78OiWmpL95xnAev2iS58NIjt3qKFEwQKjzroO8WS4Nhu
8QPO9hH1skyXkh7Xaik6rgkPjRtwF8WhboE+fWPdkCq7XdiyQdafoWO+Oiv5uETQ5gbrjA2RUAtR
z5t6NPDKHXPM4MwEkVJnf297i83QZj0bQgUHXk4iK9bcHeR/dM+I6RKKogJjY1fR1VhufKSmhEHB
pbue037tnPMOqVkSEdh07f5bzWFeVNziAUR66KOo689gsKqrkTXmiPY677acmPtU21hVS26538kk
q/H2F5dRT9so32jffbO7myJFHeQuTjh4blZUi6V7ohT2b2ZBkEiuWjvOAwTkfTW+cWs6Y7RfXMNi
s6qU2IuqoTXUAMaQRNyN1vJTZRJ1dKn0KD1CED9mb3wC25l3nXhPk/E0H/C3F6BCS81zZet6Yj56
ppk3v+LT+jKOxA0GHYtp+MONCR+bP8BSBVK+NvJiCAhBZZAvwvHBoYkeSKQ6Zfxby2Y6KQad8NjK
AQybq+sNDX2FMlYwJg8cF/pF2OtSP3j/n3dy4M3DClC5HfRX04lHTY3LhpeVX2TrvDAOTJ7u2ZVz
5QuWxveipWr1eSpQ6BJnz+UkmeCkkHDE/0nVynfGRSl18GdRuA/sjDI0nmB+HtdXT2SuzKwls5F8
KD2r10hJkauaxOjO4HJRqkr2ADYhp2F4VvPI+EiQwomJRBleVuUfltbz1sEpoGN60Eth0yIxGWaM
lItG54KMyzq3FDB8XjwlXX+8v71+h5J0Fw1EMbYP1qYrwSOtalpPfW1JpH98XuxsUo+IKDpstZbV
V7jjhC9HcizEnRaLHYoJMrhi6sA7KOdGwKaHF6i4nx6IekiXSwOglldma0sK+SNmUQ3MYb0CVnGe
tv8Fbm+fbDzmueaEpRif7y0NZsU7lKiR/bZO4pSTrIc9oBhSUcnRck+jfDVyC0dZIUqh/jvGlScd
aKwEpZO97AoOMvXhgqSmZ0hzUQgUbE6eW//ZDAPQuon2P8E8yJO6Vj54XDOqYL1RY4chCybudkCe
Ksbj44XEc9ZSdBQux9KL+CFto4NnyomTQJstZdAZXWe3viru5XBllrsFGkDSFtUsH6X50KusqWXl
IgqMMeSF8c16T/B7RJVxhcLpG+cWNrpinZwzvqETXMc6TzmSnDYaQ+iSksiVas1U6fWuCsV9motV
XlQxyynN4SkU0TjDRW68NDJ9+W93EtCBUVe0bJ+nLyxGe81jhhz9iq0Hg5oh08OopUu/8O+3RvUE
V42iKOlAmhtgRT2c1NfxhixgVjFg33n5ji2Rt74MmPFKrm6FgeCSxyD8Z4lYGwljX7RLqIAXUBhN
gFWPQEVuYEPHdNWNeAO4SXK2gVH6niRBfa3tfW6et1tmExFDOh6+lTkUzEnLJuMsMi1QQRkXBjNh
niVev2Fzlt3NuxkU43jnF4E/Ggo4ozJRjJtjAg+vx4rbO55iy+aFnTF7rj1p5uU7r++mog++lqpk
V8NiZVocuNSkOA3ceswyzwHa/zt2F+Wq/Jxh5hgYWAQmEYb0Cg/hEetDonJmP8CbsTE2yc99AUH7
P/LLXxtla2rxAsZbNGwPPmLfFXz7G2voPzXikj+uIYnLddHON4uaeYVQQ43drEwRAW15ItG70pTv
OEMYVqSF6gN7H7Jz34mEqOPWwsVcAVlL7/sZ3B9KzMA+eiD7eGEZcfjEhmxT/C0j3FvNn3iv3bI1
thMJWjqOilHXA9AA6RSiTjCwBoJdQ/N5bCQnv+dHe/U5E6HkiwJnEbLNzSo4s2o6kgZQrtVfL1r1
djUcxRm1O1l+dtegkfdcq3yN4TXkeD2Ytd/wQNbGmGIKWxHk8G11HmpFI8FUohkCJAopTsfROqLk
8P38krO+I08WlHb/8qHwR8Lqvin+3atVRRp5Z6SbEQL7rry2OZoYv6UuRAI41g6R87r8WUqIhpYo
uSOTpkg+QEb2lxwdOVP8+gki154S5tb6GWsHgFOaZWoWyUw8U2Xg/4rH4GeaaQZIWYMFW9sG29E1
vgpeAHbFDXPSAvgKYLm5QxyzsaLzLQTzyRYCxLdS11ExzY+TmCUxN2/+F+YwvPcO8tgb/zU35SIy
vJYFDA6BmIfbAUnREyph73ay88+evsUZCzirH7D8MXLpBPLRPhPwmb8GmMflvra2cJApZJbq3qjz
9+eTjAEiX6TeiyOm6mBTwuHetZe0GRfKQJBXIFAVEuPQaV/aTuDGgbuOfKgMPyQ3dgY6FFJzDv1V
p3YPBA7AB2WwmC7Rw+noko6IIsgwA3TBEgC8ryTqR7UVXwcXlDqlH4FpWAV3hsBn4kjVxkCdsJx3
ssHaXvzOdnF4VgydvEImLsh3gKfAxI5TSxsPth4ZeJyJbSXH1AyHGc8vsvayFK6zoV69tmzLj8cD
Qq3O07ZzMjq91/M28eEo4tNi4x9woUznjHcSbpq1u6Coqj8sxCkGFsOTMu1YCBuCSzvmjBOUkse8
/nV1UPDQb1UP69HjM6C6MP1WgjCokyurPrSuSNyFAfZYuAPZbEkIA7XJhjZ/ONJjfbPmBll9FMfP
90lX/8fJYsRsvLbuAtmTXbRpljHU2MfMn10MQznRTgJzhacl9BwJ82Q5AI138TURwTd5Y9wZlu72
GWdU52Cx8l2wYYWGbXDbIkO3LZEGJvNCYb+QT6s8rbT4UYuTNXrQj0j0pbJ7YZYE0ts6EbIDixUP
0Ih3S3H0BdjYe7Iv/yHBnucvLshYKzkXeM3VHiw9VlP5/ztdczFebjnB6ckA5UaOU6IM6AkjvAaF
iPvltyMgHD9/BCmqg94caV5z0hOSgIdO5K+7VCCYC/IjOpuh062ONNtaXt7CWgTAQJlmcvBSoU1N
sYeDiKHJA541me23ua4SM8ugHns4uYLKCfJMVardAcV3X7IgF8NtgLZ4L6vI/mnvRqEbL8BZQQAh
h/zgjwG7P8fN40eCL0shYWpTuvrfWE7+U5FQ4Ptfr/jeFRr2J+m6c8LKzmM6rWOhu2epC/DIev2+
OVubCK5e0uV/6Yc61nxamo7hVmkjb0LKvhJ3Fp9APz68Y4RyOs3sam4/Qp7uG1q0pxOZnwta8Rtq
aQ8FUvMbL8iXtWphNscpG7AGBsszISw4dMqawew++Z4XOztvSROc6DwFHJ8dhCCvY0nlcD1Om5ST
yP4Vv7MKx1bD2HuhZtF6lu19j++AJLMIvMpyavf0dQOLI2dikCeEEPxFzh+wQVHGqBdShuwuPkQ5
CwYgXbdb2S9LwFxBIY4nZmGKlEr1jfvZoegMaj46GyYEQNyQzRfY/UwL8bUbtOKR42Zo/vRxRUDU
v7Px9VEX28TQvMl3f8h2A2oobvXt7W8iFVV0/7qUztijKTgkgVfqjoG1IDlwtw/lrwc0+XV279fw
LPpBFHd7v0qQ42zis+5zSGb0b9TmqT0eo1K2wKbC3OK9dJbeXqV2m5p/BPYnF2Y0ML4rKmnqnKDU
2kMLQSCAZ/BjAoIHIvxQo6Di0DLsSCLqvu8X83aGvaA0le93VsJbr136/fRaxaeD9Irq8XpO9Cka
lHyjYmwvRFOFAvQSf325iK6nr/jMJ+0vvFGNMiW7l5jHIxmrc9Q/ARHzzen4DvJloiobOrIPUsUw
kNWAwzkKrNHixIIk9mUcPX0pAUIluHZ1ZQ/YzSqEIIY1DVAZ8SEWJ7nsY7fOeVleQXs0LJPm2klU
fPL8vQxcaN6FXU9bwvECsPGT5XojtfUdZ3FNSNPOdyAk2dX0N+RxlIlfDHFl9KQ00P+whcAO8+lb
zgZQQCd9i7dqy8HTgTP1idhcYRwQc5BZCaZViMA6VKSdNwvyM0chUnOgkTZ89VVq0rtdrNCRPWbQ
KQOvREBUOTlVcI3Wy46JS6BdHUpFG86JlFEqIEfvjVa+PwDPab7q+JHGADR62pp66mXa0qLaWJIZ
WkBk40qL2ioGb5VMmSmFLguSLrlMEwtKBU6xcNUSaYFLdcnk1YD/vs8Cj3aDqofRZbFi32FOsymo
vAFEcvcrlYXtcoSIs7aA1eSDHX7HjTBM1bLif7rBOrvqHv1+29uaXFsBtS9p1En+JN0kKvbmZn3y
MqUhippt7q+ca10UO07GEpOVc8RhRQaPkYew6T0t3Z0tKDkfrYo4bgVDetsnbEuDvk69N6UO8Hhn
P3NFWIKY/kh/LrrSgIp32rv7N2LoDJYXVjmBEBxjGy42/ccultTkltibGou5v0lwyL0fQCojC/Ha
kyNzht+MFjt50ChV172J4wq0NtQq3oxEBqGTYxfy7fyXimlcjful5RDrZ+0kR7OiNPPbrGg4YWWp
dCoGRPRDin6ZideFWZFvcZkfeggXVDd7gAXwJ9aSl+tcc5msiFxp5rkmAD9GK5HmuBKfkMn3oHWv
zH06fypEclhr31FagoIcQax4VHf6XnJoSGflaNtqXlvItZfpKlYSTOJ5Ng135yx9rPrCl1Ccb2w8
AJ1he/sEHaFWSVQn06Gyy+097aojVFfq+8dJNKja1fMC+XKfHud6YFnOefhqhZzVbTOX1RVH2VWT
ftVA3/+OoD9Dhhmh+HG+HUQdIaANvRan8sCg88zNyvCQSZ6AR+XyMWp9xLcvfjHjvmFqNRJNXXRV
whvHz1etuMo/TJpjj+0SRD0gxVgq9jdVCdXk6BxIboOkbQQ5cX6l1iofnjYzGDQ7NwP+RbG74lcx
14VwdFLdK/JgTrmUbH9D5apheXbDeLFQcXaikTU1SwKCHKIT9lsC3xJb2OEi39KnDAu2BhWieary
lE0tDFMQSCib187Dwl9V/Gv0Z5qdn4YjtHmBgrmO1/EqN3h4+OwR0xT04M8t+2/HojcFsaEuavzz
krP3z0gEtMS4djeiGEt+GClnWx7Db3NyQ+MnfSxcAYv0BDTZ1yyAP6/bIrGonaLnXBkuwyQBqzaW
xECU5twsXDlYN25I1bLAeCo5O5MtRkw8yiKJRjb+XXbsh06mimyzKvp2wbwqiNqKClwiHMqxtd5B
quw87RK8BUTuml2U+lkrBwDI6Vjq62RNC4FXnRSc9zGL+ioIsC42p98YzehE7YpRZgAliw/eJA/j
4cXb9PojclJJ8jPaJAxnNRFXAzMP7jmH2AxuPaEP/da5QExmDV/MIRXxv1GLrYNRY4u7xhUDMb+P
paggtbqDtbctHOarnXkZhXDwFTyZc7pqn9Suj0gK7cBKNF1WsVfHOj9JTSE+Nb14Yi3sGwU+x2sJ
4q4kOmKzMCNT1OTCrmjAJFQCjFAdCHVGuCb6R97y+6viP4qRPbVuRS5D/WVFxy7rTq5P9oUNiSgw
gGm1MHC60NKBCJ3bgjyW4cBe5XCY1j5bXsjWH0EnZmfNXKfaEqOXvO4x4E6uOaUVk33Wwu2fZuNl
gjQ2PIgb1OG5ga31KDLTot6AUGfWZ2cS0W0aAKXps5ukVapDTXDLBRvu1bOrijGdtLcdDhHpB+xX
pJzoD6qUi7KG6CIDUPYfno6te0HQyfnELDIAGBt9PZFmeyoLmuHlZ1kmSfEmWY+xMkj9nxACjxFf
9CWCbd9rpgkoTwfL9WVnNNku6jZLNgyiAwkibDamRRSpX6DbS5oOUtYggpM5jnKPOBnBjsPZKEkV
BrKnim1UUN/jHQ3RWZGl3etUNHn8kuVsIJfC8UuYCLZO/O4Dze+LhkebSSfXesh7VDntsreF0Sa2
2O/PEIPi5RU3Appqk2XpMBaAPXMpK5KHN2679VMKP0va/OddOij/BBRTXLcb9DiyFP3brDwgz6AS
cy8KyK5bYvOFS3viDVasbZWRJVWPx88+NKn9upeE0MwqqitKnhKFZJyRJxAWGuCZz2lg/Gyob6Lt
RuH5XUkNBBfTRIAw3BqL5RF+MCWdtvlVwOIrzLNMrAtL0V3BGVgYlzLNc0h+zbMljyq9gYWg+Qln
+RM/EYs6mtFoAOESKKHyYvD563q7QpiDVglG2oqqKAWUV7Ahc+XUITSfyUNWKhSfWlN3XYilHcf0
yGXg3jKw9zhsU3MjGkhWyDc2zMw4Dr7GyBcNAI9nqfUbzhN0UyPDB9kg0EHn/OyuYJ2UAtihXGhO
Hm9NNfO2Mcp5DtQf3zd8Sbu4WW4vHPdY7xJinrRiBItevLTt2VTkcxfGeFwZuitwhzPihg+yR2p1
YRUFW/ud+R7a/szKjiEO6ZSc2z2uVIK2zfG64VOVxWB3MOclfbgHKBa8s1Fm1Sz+DU2ukZu8oSYV
zZAVBu3J5Q4Pw20Exjs8wXgbjfeWleAVMlItwQyJn/BJD2vUM5WX1Rf/67i1WQy57n6Fjt4Qf3tG
v8si2GM9GRbbNEqlwvUgMyoodzDY5xxVR86+8G3EAZ2DMx2zY2NpLEfCCCVzBn5jnauFoxyuXEtD
t5pdehpIgUaLLcCUblju8ZfCEm/ff/jn5CwG+mJa9EuwmFT3cY0u7FSEQ29YJ+8nlMqTQxkcvJh/
DEfk2N7bcOWgfpyBZEPm8MpLcadjmW7LMtncKo5JKhfOlHMevT6OGz/aWrfBvEq4EBpgdgU0bjxh
HHWE1NUusKfjl091f4MM79QhbwVDfKuKbpd20lgueQjSfMB0oUEG8bKSwy0S9OEVn0SHRqWolSoK
PKNc5WW74pz7MhgvPsSdGY0/CT4iUOGt4HoRTrX7HZQB/CLONY2FionQiEl6O7nk+WjbX4csgA3b
yaV7LdR/cN05v4cjCmsIqz3ktFbkjt1qSMmqyL7Rv1IDkrUg3MiwovRyyo/mPd5E5wwkUizaaMVh
uX/NS0hP2XK7zcH8nzs5ziYiU5SMIesLeejRjmjVjGo4lvMX4m5H1gQhW2oloY7CsHtqULdbyRBQ
0/sOyzIExc2+CWyrx7MJA15mYeaVUjQY7R+ofnP7mAn/mQ9Hvtcwm9caLYJqNkl6IhRNQfZZWD7a
Qw9yDz2vbS0gYAlJmWu2UOvThgtCcawZXul22rD7McqhTgTu4ui8qgCpGSQsKxUv+eFaGfumRhgc
sA0n3GjwXjIMNISp+VEk7pKHIlri3fxEExycGdmXIYIDIu9KM/dKojHnYmkIK4WU6wbSD7elX2Oc
JSGcSIzXo5zpwbPhisGNyq4ETuz8FTP7RGoYFjlZ7SXc6UdGzfS4UWmTsyGgAwk6FU2wM+hZ2SMc
knao5SaSFysxVAIQyW/E06zVj3SKzziVrP0uW4xo1um1xfJWw4M6b3/9fcI0mmvys8v2rTRJ1rRA
aJpqSQhiltHaWfeiSSBW+t2QN8S8Sbsc6xD/7FVQsnQVzFvJ2aptgZuz5mXUlVc57Czu7bFhjqQs
9tyPjbusj8CABOulbb4TLS2Yb3ZqtpcreE4/SWSAXJa07ygiqt3JwoR1LW371nNjMpmQ2OsAJJbW
xSBdS5euUObAHnARCWIkcErSAX7TJNYXScC3paNshF80TVPvBcQAPDMlw6vFfczFLEz9HyqKbyBY
0wq/BpP+p6yJyYESJawbvEFz61u/1gS40SKY+oMXScUMijWF1ywwMeZOU8sOEiMc5pMUli2lntxH
MSWyZ3a6Is5+nssgwZ5qOGoDuFZYu35MRq8zW1nIaWThNeWT50/LIMEqCbw9zUBDbDxrVPo8JO2U
fdgZJEzxG613H4zBj0S7K1iYCYy6W8tBhrqP4RVTnkvJ7SLOkRHCd5abJmnNn5L79IZy6QHix+y/
AbPJxW4crydsoXtDq0yQjENrJYzAuiuxK545Uu8P8TiM8MDlbe2cwGRbk16g1U3nsTweFr1UzpHB
eCmHcOmQQP6WjazbMde3BBnc8kgtJkFsCXljCtk8Ch7xEhkbtJ4Mb8oMgOzQQLw+MgDQGKhRXNdF
yifh1NWWyq962h1WtZp+vONTqPxq5N44kKFoZ182oDGN1hKXQVBJjub0tneqnqTcExnzBoNlhhZz
DBLCzWSEVeovg54HzOkmGXO+8XnZ5SB+UPAf6x9z7/4/B4OmniPLW5Xo5mMRoN8sCtnzBdBCXrhS
RttHh/a0ZRfaJi33Rv60UQjtHdyHAB+CRtk7Bonsz9tSn+wvzN712UfQLVZ506TgTwu/0oKgakuP
Bi/8b75JH/YRd0Ur+4nSHIHZkMTE7cqp8bb9wbaVZGcpKZ+V/AhdNUvwFDsdpz5G2ttoS6ITDrTo
qrrrkTzkOQgn7W56UAfV1wdC23ivF4yPQyIczXUZ0oyeBPce2r4kqCDBwVqdvtOfStFcajRe5Wb1
2xAZQEj74h0kCTCFrVSqFx/hLp4yhu3DbCq1bWuixNM2JOJPjynzwoQK6WkGdGSvE7ZH11nCX52s
YDz2+edGkydrQXZbLpHRqvyQ44YQtjgaFiQ3zyDPvdBkHwTqdmnCU72YEa0Lnxzat6Sc5mgxkayc
biz/OHkVKaMKS6o3tBrtMvpReprG+4u87pXIxo4je+Icox086wruQ0gaAi8vYx9RVrBAfeyadAF7
NoP0dvwILM4O9sKokuWpGs5KBiHQTzfpUIkoB6kZGL1I+0eW8o6iZqmQ+UgJt5eorz5fJty97KdN
4edIvBIXEDhiXoFD86nufATmwB8adMkTOyul0tcos+w5cf7HFbMymaJWUtVI53d3Bubxl5ouIZaS
bFjDBp0V57KZQMk9Mpit7UfeUTPbaZHFF3/88aR9afsd/v67+Rws63l+68uoutXnkKPnHljiggSc
5bq10BYbUjqqgnpIjxtc4VxfkQlDvH8Dae4qtQOe1huSQVDOip7nTmJhVgSC/6QBP/WQ5wO4zeCA
+k3pf0Bcd4UhUzPsjIZwHali3jSnSd74KH1SBKVy7E2bCT2g+/1c7fqhviqhUcA2rdukh6emLFCM
K00iCqHlCk2g8H1lz4UBoyFeQBxLV9sBU9J+fuU90kD14Bf9DufFnY8xkIyOTIocQ8yIpaeHezbo
m45aQ3pmSXSqKZINvloIpiRu2V6DAib6Y+RAeC45L5ZCv4/uEKkpU9c4E5CuVX+m0rHFQV9861Hh
fyTLbYC5Zac9XDMoc4BGbZvn4NCez6itAyeOLfjRsX3nkBFIvfKucVYqfzMDZc16SgqBmj2WxmVf
cBbKYUB8FdP7zPJKVx2kB7MIrg+5eCDFvcu0L/uVmhBfbIhZxInp6Yt8+qA/DKsivVbjpDyEYAt/
0vUwaG4bHjZ5gwjEHAEjXbN9i80kOsfi/+5yt3U1yNUxZfc6d4rL8jQ+7JkHaO5Aki9XQeB38080
rxbL2MVXxi06+tO0vDNQ5/Hx4jsGRrFQ2SwxDxYejwiONKAGEGyyfgwI9iS3Rn5TJR+PGndl74mH
mWPlOyB3UloHw7Rnbx6t1Nkut/jegkez7eYH1WLqGbNaRbVu0ymOepxKfsePhYGsayuzDlpa/OEv
aUtR1iXXnuxVsdk5KNL0nukjMj2KDC6Gis0MC2HmFoshoaDVhufMRZbhLXwQJSQwBK3+TkEMOgbN
Ep4s212jCY0kjKcg/1Lc+t5rVEX25MzrGgp/giCVOEi/jLgyKiLsJZYrmbQA6oQmMdxTnh7D9pZX
/8vgGwjouD712YL3nqGW6VtM/sevfTJaUkCVEkY/Yw8HWA+Ib11KJBJijOtw2/g/PpC1NZPmtmrG
o8pYo/IpbtCCH/Lm+Wyih4sv+RxPSZH1eKFHq7xO1m6BK0AmPP7OLAtwqBLKGoF18YRG41+MQJ1d
pekDPw9FZx0rPncLpHtItML//1buORWzTqVKSJjMEDZTkfwAfUJ/jC2+u1TuLMQ6+ZxEf8h6LCvC
QOYg1zyqTX4V0EO1Mg8UB1hUi9+doyJCmwkStEevwRfXlvwRntg9a/MAcq0+5ptG4vWNpUwasjng
O1bmjX0Na3p5jK70/2226M6Bzwyj7UucTShdn/pIM+tJXI4JktFKduhdpPTeiRgGlcoory6mkPTK
KQ0L84sWVSHkY4vlLiwxRvwBX/rKj9UeovPlxcpaz5wFBsoJ0A9uPorz291AIn3mTdaUEI319ngU
tbbPcRqd1zccEdc58tSBwgxpa8ZTBmVUC/v76sRcL7a7uAhi7NnaGY/W9CAoujXwCbyAsrWor10R
OhLzyVBqER9vQ6mKWxeidboBk4J/vRszPogaiF+Gdfr5LunTA89YEyJbYSQHmuaJcqEEyvb1FcJO
gP4o1fxYUpCnDkF5U/V0j0/Ke7ppISE8byIPZhsdwbkR8xYhxtWwc1TM8XKe1Kta1xiwu67W7qXA
WIjNPLI3jz9a2xOy5p7xkqrVI/0SwGJQC0R4C+GLs5bfPtFtDceEeb1AgQI0UPMn7tFgk868eYyc
IsAmPlFljSuscwXFv38VGrZpVS3oqlF3AeVdjNe/2BsFYWmZx7ElUOV2WepQW64OkPfIpmidHDz2
X3csrH5Az3NRGXrtglw+Q/LOvqmbdQ3E3STFGnheIrI1juEcMeCZEG99eSEPZNyBm1O3Yeqyy2Sm
8xKytdln+FheBn8n/5KbKUTtP8uptAs8Hm80soXWbu/rQ7xilW0f+eMAd4v6LooZ1umPUUBpwnJj
Q9leX+6gsi66k3oZcDxomxfEmZuXa32sJsI8saYHjJF9PizhnCSPVYVIyDZOOI0K44V7fGoI+txz
GTkUy4oAMcrF+iUEsN9xRam15KVt1cwAU9AXhOPyRlRzWDu2thOlqX9SZlyU5uN4DItcglPY0jvV
MdbSio/z67xMR/5XTkQryzSd95O3VOr4L/yvShfcVzz5eBrNSnE1zgcGIpUWu54lB0GCaRUx/197
LKSF3MOckHqbm9HdZqZY9GctacmaZ5qwNHNVSPLHr82hom/s0BoHGKV2V0vJbN0dkiAGLC8csHR2
xLKzfFIgWDpmlF5y+UfWiEeZ8fVZTi94xWSEaQSOlx4HQ0ewKGmPGKN02+pOOvKA/NE62n4Ksh3q
0nxp7jcmKCwN0Gn3IeYMxRbIVTqIoe3UJsCtNYzOrNnkK/b9vfF/+vjC1eJANSAq7KYU6TT6+Xp+
Z5hvThaQ+t16S2MRUymjzyYhs8gJ02aT+h4LnTrISmARCIMWv8yCuPjMvUAt1G5U54SOpuLV10Rz
ddQsFbskTQmQ1wqJIcrLaRccVTR8MDVTnH6kqYQS6uxNoYiYeg1LgE153bhGMixBQ/KUkWdqzyu5
lNytfU5wDYmLBWZZo3WzN/t3UPNmJzu/IKLTvZkDMT7HtSEgmcobv9KN33dYvHbPTcQB/S+7yxvi
/MMDbkrL6NPTgrMaKhv/yi4HVPyxoG7mYT6zrzgbsEM6l0jaBe763lvUpOAhRJFPDpLV0Xnazky5
kT3sTqJBUxLJ3rp7LZd7H3mp5xNHGs161YHS+gQ8Bz9rgokH8q4nH1cT8ZEjs/a7EIf+6SXh8Bl3
HMvevBzuFAWE3lwAUG5WamgufZkDP9qsekNOOrKqmDWXvv1/zm1k4VtK35Vtvb6lXiYZoIMTwTwB
uOoSLyldTMFZQzktN9t72Ai0Rd5iP9G7LU9THF2NNx3acOWGk7IP+uIwqP+XmF9qMuMjDylj8hAV
bbndKZomC/n0ChmaqLpS0BUiciUhd5PZ0wWkcQkIIwMqLBzthoS+um8KNYoPkDIIRUNFNCNsu4/w
ZEFYZ9quBnfzHp2vgXw6FLJmIT4a0iANrVyBa4gBconk0Nvs4/WInxZh9aCjRfMgFG9BoYJ77jLi
bAV+cnlmKrQVvZgHW//UYu2AmIIAb3JBkC13PftEsn9Zmvm/6eGJLNPD2R5mbkcPkypkFWNw4WTT
XDmrOnfEBpFHI+RY28Rps8SACvV93paGY9sx4X4R0QzF1SCrtCp1jzxOYXkbEEneA93W5AezvEa5
pkiVBPq+3eNGYSfmTBdUSt/sFi13IUCGfiptPbXdUiAfP9Q2QT+VBNlFGKxvH69zvQaGXo7okRxF
xg/H1EuNe+9GICGVynMUsGaGnmHc8TuxRdweUm1Y4q9oOqAb7Xlx6L1sBxw1t0JR++w2R/gQhPqI
xqvgL2a1x2nnNQ24jh9h7kP72KLwGn1zE5KQde1vbwCwH/UCtlObmprZWZIVl1l9lb/aE/lV8wh3
ukwY9mJWv0U8eoacx/ge5pZWTrXa+5aSlI/FWEvtUasS7GlFIFd1SA2iqp7pKGV0+SogK00YEPfN
zyd6O4/Sq7yClyZPdkTwVVp5qO6p4T6mDlBzwktN/IYwnby1wtLH5s0/Fnvn1NoF2l6zYw2iiuVb
MlGTj+iuFLvuSYXHS5obWp7znjpj3gzv8Wkz04gacjJPjuu5PUzOdyCC+IBxjMvvnnezJaIwXOOk
cRBE4G0E7qZqDiDH86sc3OmLiLpq0sexYNY/0BsXx1/vuk867sDEgXwXbM0sI4QKxntJCAWbsX4H
7EVdNdowREmeCnLfL90VWz+BmlEnCk02dOLvkd7wt8CYpFzkLn996IbPAaIwZ7SjEA8SIHOzOb6d
ucFYICx1b8zvoqqmaspWLyj2CjYbds9VhmIv/JZKwNhvnhcvU5zxfXjtXegHYwPf4Oh+s70+64rJ
c1k7T4KFcSxIPKlwVDnj+FlOxphdPA0YBX1fflalOHpF7D3OS1JDHeYQBKORm3MQxeb7OIs0lZZs
zSJ/Wz6k8gJagQeI1k/qz/GzzUGiRi0G6EfgTq9/ZDrqq3mLuq+TOBm23f5BuGJAoqzhaL9hRqk6
KohsYKFXY/2wdMdu/KWJWnkkBM9nrbQzZ9L2LJlART2pbInJx35cQSNLUFlmXtLBkCna6zA+iepl
NUBGQzhw5DNSep3h7g5GZBNNGhhqzPtBmOFxSERt9WyNkc/D/NU02ofxKjRvsGAMqdYKVLQp2r8q
8xUPowTa4CU7VptZcjtdNSiwrKhnxv67gJwJa1hHBvzF1ukOLtoYh263rK5Bo2T/I/n9YOW4/YcU
7sDggLfv6PSr7Sxma3FXTQCCup0k399JlRQ90MeENXNbatsfBRMOD9t4TsIfSig+l1+i/9Of99+B
lvbwr4YyvuEbBUkcNazapr7jXZuWIP9Kyt7okRKtYVunwkTaNRvclgYj8OBJIXaibKipBEwyCQLv
jClexpd5pWAH7Wi9B5EpeE9pX6ThCgjxJ6mwnc5wA9cjBmCZQshxPeYaN7VNrsytP1IHEl4kuJwb
TbO+ymMcfVjv6ubD5PbRrfcBHuozhyv5/IMKX98RTyxZL2VYv1a0jlSYA6iOQD1nwPT+o14y60RI
J/qf6l/Ls7DHP8xHcq7F2PsDNsxQSA/+u3CfDVLldcE1z6yAtIZAjS59NdH6fdtTmHXxU3X0W4S1
uBvJSZAoK3D/BHp3HLDgoCaFKhu3FASDNvGOQcv9M95X8k2SlGonymIHba1K5kGLMRr/XyxL/OIJ
hrEV8HYvm7qu6jJepB05+8BzXWOsB5bgf2ScOZjHV1eNMCeRNZiAVS+Km6pCaZ8lWSZtYSpux6Ok
7dh23GT2er5hIF7SBF7L79oKxOU4o71KlbqMVvIQ//hNMvVb3J28C5wU1GJFZLkxXLOyivl7OC1j
ImvAxnE6qYVS6PPmnIKcGZnKbOQWJ/A0Fic6daSpkIC09GChxYeLaCjhY/IydAXCrEDGNGYdQBD3
9SVAXVgeMnZ8HK+7lEh9TEHm4z52AItQXO2817G+XIzijB6rfCJYG4DoEu+XWBbrS7pmTlx+pPpN
wrPic6ZQBZVAwcWkjUTIR89AydGAkXUR8cPhFktyJN6ckQPCHk4vm6GWmX5FsPB5HQ9MQiFJBSpK
kYb2YTjdGxHjKNjbav8QyQm5ap+E9u+aqLjzDFuDbHfAEkLZrwI4yfZJrksbsodBBXUxYmnDH6KH
iqxTCkgSNyqYC34Wsk4YPBi1949BXQL7RLo6eUDWl993OoHlET6ouR3bRyQHz0TPuQf2kXoHgoYw
I3NLZAHkV4Q30+rSeauntS9XNhkosPZHtLayFGPQ7l1OWRiIFLzN2cEjo9rjDVU0/sgI3Mx7+hcA
TNnOSYFc6DqtWQvarKXTm+y+1JJXKLvQNEpfxhswVGudkKIenyjyOKLmsqGs9cNHalVrsBjqmS7f
ZuvtCI/cYITzcUpnD8lbNVkJMxibphISl2YDm3st17r5Jc9iiky5QKnY8UbzC5GEjPmU7omiU8FW
6yJOtvYmpGE8qSIdg4pwcLJ2Nq77mvWDRsDXjpKEUFZAys0icIBH3Z5lihyvOU4P2KAJF1dqKRTo
UcGnxKUYYYBFEsI2pjxD6Sf03UX/FwEkaK2g1QajBuhTXFvY+HfpFsbuPtj3pCzhuRP9yy91TLdF
u7iyaoM0GbktcVMmThmJM+iUcTagDwZr3A2pTCUad1lQmvdULtunudzsUukJ+8cpz8GDSkmrSGqJ
l4CJMoNFY+WVK5Sggy9KP1r1LwrNxxBy7eFU6OGEqZCToAk3T66I7S+LHBE25k4bblWhpOsnNRbi
LcsfpAbJkakTcCCfilvUe/yGTjCt83dABTmZbH2/POT82i4h9/GuE8DJLcGSu91DNXTadRuOSp2b
o0wR0sRE/Kgt+0W45RM0bn4J4wfadiyihHH9fV48lU4gRhPxSY4rEWvL+oiAhZECvvoKjdcOENBl
rf6F9H0mu+UzWiV2EX/0Ow50SdqjLKBiSQKFopyAaSTY78jL+myJ/Ow9TMNykWN4trWmzn9CxuVa
We7rYeOqykwjchnKM42rWDghkXuerdgAF2efJ/D85hiQ84mYg9PQXWkDRwWX6cFoL8eqw4qCxFRD
yvhuxeuHaBQGB0OreVV6lZkDiPpAPWuXMlq3RbpH8xVOkJckSaoNVjL4kDVqHtAgtESxg9xu6Fup
fOYdBT2D28e1AXYotWw9fZMMnhAm8KHlOCsxs7WGsi1VbGcgml9eaKov+xB+awxYvbA6G8c6NCzX
mmGR7aVDzSK7GRp6CDxPnDxw/3vU4DwOHnCtrgyjiJe52Qx5F3pubZR5wm8cAcSTSMLNdCqwqr3K
6rSQFayXVKp2bbTsn9WX0aE7wIhh8efZj57Z7k4Bu1h2fcaFvjRajzm5960oUYyVRyqY0i16mPkc
yShlyAD87xIEmLzKeBsXEvtAsN+lKNOd8+y2QpYM4YLA4L6DL2K/YNG0D7leDdWh6CIBKm9rOCKv
RxvISTm3/VpuKCXQLP9NXKUcSTZ5uv666ygOV29pvLrHc6De99BDlLwrO3FeiTurXAw3aixnZgM3
eIH1nqjYPx3ytAXom3mQkcZITfOk+95Wmm75NTAOSdQodZyKKDolUQeT/Tx3h+0rytTZ9fJffqbP
g7bCZYE0axSg+5MqGdPut5otUdOAcu9NpbXEN7TFMWf/1VorH6+wKmQqdmDni5tMAWLrSxVI/XxW
ULjMK2eoQcyi7JWVGo72eQZ5040FlR52l0fH66etvKge78NSSV4p1jYEBjHeFDiDBFeKlLjrkuPk
AgqTETibPI77sFGVpv5W2lOUR3WryHU6QIje8MHWAiWY3fQ0WwHueWouEsDoLvuIRN6VNfZC4/0q
qBHE8JQ+hDLhWdxGx7DVeGBNcO3tx/LhJJJkkZ9yUrFngrX1fiNEfzq7hb1u4CHZ4ywymwFAKB7F
TeRnvYTYLZt2lQOwMrSokQaodr0BPnA0lN1GiPMMFaWzdoUgaQ+upAe9UJa4CkOUG9fjDth8pCNK
e9L+o0wQ/yVdQXTYsZhlJbNOhEmTYc2LKj4EcJ8twpVtxsZV1zXPTNdR4B3UUqj57vlG5p+XxHCW
b1p44eOopW4T+0w0ql3y7gTdrUhCNF84+JUJDRv3G+Pnjt94Sf1SYxw2ihKtGdqyzr+iI3s7vzr2
ddnsRLoq/AxEdRvxpEJUiuRyU9Ghllfjhm7XOY/m9DOZKrJz04imNuQUfZr8HIV7CJU8uHBOFx/H
jK9O662rA7jquXwxTt3HcHz5aNag6YF3jnzc82UTuiupm4l/5sXRG0pwla76DzZByP/VDNu466GC
ix/htvetp0s3eP6Pu2Utahwv1pAU7hhOvGiJBy1dlmnCdhZ6hS/gWayLIYsWs6sha/Q1hMhzLwj1
kq6xrBEZfcvxGmFj+dJdb09jbaABAd3Y0+wK4+LKqHeZscVtNluh0HvrMsgDoxqwg87u3KGTEiK6
Z2z5Fdc7BJlQYebPqtjWAF32GcB4cAWmjgJRW5TXvD4+UjDO8UKfPjzPxor5iXzJoHGnc17lvYyB
ARMyl7bovIRBPqLG9APXUx+bI4kCVh875QI0Ims9lr66VF+l2A40L5nT5hMoueSAeoIm/u+1Jq0r
Mi/QNq20dgWFPo+F52rBB3s3TCUbeMIAFUPaxs9x10sMf/b+mx1ZpqH0R5RCjjMPC8u9IAbZKU9q
p0i6uRUeKqv3jQx8V3mQOLZtzZ4eHjRnMZPQE33legVh9GTQNQrx+W6CllLFTY4G/02fGk3r0Ffb
TgOsEzRs8O3MvtjGy7+0wXbPE8Eemjz54b3dUxBdEJP8zRLx0HzHep7qTHAVm8YhqjWLG1I2x8L4
2aWznqWQrvJ+z19NUXxqIxmdERiosUr1PkEVn9p2vhxcFzUWdUJYPSJYbUEATo+AX4GJXQujPrLg
5B+h6hlpvaUs+0y8IG/uEZcF+yxXLT863xgMuis4F73xFdTOc9Kt0RMPWFwhw5R+AYR5xF6dKlFI
ni3c7pboJ4ipZ3jwkRMPJTQnZdE2Hn+GAvfxBRjca1uwlOWrzhD8kdqMi9IcSMOT6mC1vgcmfbHx
hgWPS5X+4c/QoYWaFc/hZyYJpmQ7F3x/bJ6lb1TbKgN36ybIEtwapeG4Lq5cSobhlkVtQzUgyPDg
a39B1+4Hr/7ER4l/Er1/BQtMeDFpEAJHXYxRgbbX3vBXTHyGEo5JUzlA+l1Az0qYpyywU1fg8hfN
aVtuNFZDTu0aBPEKWZ++IFTFIwg8S/F7ThXtz6Jgyciy5RRcKowqcv0BtKfO9xrVnJb6aHo2037y
9wn04tE1BJWjcTyvjLQ818c65XNsOqYAQrFyF34ol7UfdOOY3M8d9elNN0aaYJwYSPuz9z6Shihf
shmXrdWvgYzLT+xZtUcr2FzV99HTakBhVBbPZwaOflUMuo8DHPj712+Wdi9cBv6XGcH5I0xfPuCo
2s3QY7NYrMJ/pacA87SgxZbWrgKmT9rP1IkMIBPo5ixNPwEtrjjw1D99R8aNCI+vo2F9Aq9iPbpD
eXE/RtJliN6+c60+2TIK0I1LyKbLvvwF71N/BJudRZMF8XLJE2RQsGFX3ZK9hDiEG7k3S+Q0K4tZ
HmrFw4K0aYTch5d1zt3FJ3Os+201TDkpwmWhqyM2qBHDpnkYGEyOgEeM686eVPlq9MaGkql1VFQ5
JP32PUW3KcnlmsUYZ7iJSHkJWCTpnomuGVxokvCR+CFf6U7ugSS76VDL5TVYI859i/ikySFmjXf4
GiOwrutC6V7GqlfFX/ugFNAva2wFsKMoFUK+ctS3UipEtzo0+sLfUm4l82UCYRw3i8fFWH1reb9N
jvc+hOAF+AxwaBuVJjfof2DULhCuNnXesIA3Vhx+L5dYhCNIlOMVlSZR9c+KBG+ELRvis33v8meF
36/tXjRj4StYFsIoOlqigBDEuMA6F2TEPw1EeZyqBi5Ma1h6535l/LLKVh4oqouYpSmzDrRK8Uam
7HghreHDzt2HW3Mv9DKjKtaDWV/rGn+UtIJ8xUduPo1YsZL3aKWegvDqerf3OnJHqsCHckUgKWK1
kaTVBJy+77tEms0ucBcuo78iVdMnFB5xxHRO7itCa66cCYgRmIv5MsyqVpNJ24e56ndsdrN0fRbm
jF/ith1wLgunA3WC7YXFSlOq7RBEC2b0k88WvnnqHetEbnfzWqm2j8MH8pfkjaqvI4zQ3lM2paq6
kBuwIa+CIgtxHKd04JoRsCQ5S+fcRtf7Khskmm4r023YuLJ9Y0qPyjaRF2zC8R12Ko/vf48UENuH
Pzueyqvqa8t+jcnlCKBO792lF7jhJhCMF67iR8u+2LdS15eUHjPFc5DvABwuhWbqXTBsIUHMUeut
vaKL0UTuvx9709UlzWFmcTX4MMNvDS3VlKQa9kUE1VWxVbR5cPgWQ13jNXZ27zHkV6F/SOYR7HNN
XsEPHIRLjwSEE+G4OU2m3e+aHFwdfEDlgiMUc+EgF1mUvE4lkyQjazDZH8HCocj28MwCMbbzaXqp
aWY9XmfHjY+/25KCRgCQPb3KAlFFdRHqFbSWRA4L2uMBzjNAoNUy1t/9y65HsBQ4uxtTSdBlNE6C
uCmjqzHwiNLgRwZpZwmldxTbCF95/lvuvO5i071mpw3ksBech0LtkNd0KD/hi99j83aG7jVPXzk/
CAAtoPwf/YsQjQYBw0Q57e9VYa1W88YIG/Ypdt+0+JKc2u1Q/zaozWSTrrJC0ACs+gUE1gi+7B+c
SmJWXnVgbr6j6rJQpiKwXI/nsY46Z70yRfkSr/HTSdUl9POhlWSGJ5MKswfgO1zP+1RXeUvM8VpL
8f9PfzHHrU7JDoO6Vq85pivsfLXXZyPfzAfAsM1/7H8fdhmEjl/VY3zol6z1DoVOgowRO0lkM1NS
QF5OSJzLPuwA9JkfrvnTi1NitPoS+sW56g5+CmEUgzZF/8HE42L2t3J+LsBiFJsHEIOWZ7vCqIiK
pOM0raRK+If8pgaJnUFB7Idw0cve0O/R0DPLSbjpBzJ4fDvkT6ejOtvIUES0bYY+96j9ihNzpq7P
4EES/L9mbXg2kCqroGgDwqTjcbkwP8OnZfPtmFBsuScGjxrm/0iUin0RkTQmP8opXRtGhecQYjqU
fD4PVzti/pYb9JmFCyncUJoADPafoMJwmiDz8VO6GOqlXNQ/NtfuI14/jL+Xmuce61D0KV8cH1Ky
qXA1Nrp7RBxI2QQXcQS5ielmH0JBmpxjt00sHYdCwQi5qr9sIt75d+CnKEI/SjYqKgRq8sVGR0W/
hNsnCSzcIN53gJuNNdkFqCv4a61PpFK+NUfi18S+/fxpHCFmo3N70P50jgFpST1BMg8FVx1w2MiH
vZi1gtcD1oss5AVaQSSi8D5/eXmGvgm1Wj8HyT6F2NX08BpVDL3dyCYsXSrzCEnwUkKI+LO2G6hE
sRuD//gwKvXK8xK+8W8/EEU25CBPjq0WsrR4V3gxJAeyE7M4hdytOyCi/nHrjPbSJczQv3IMn1Gr
VUWfN4sBaD0kL459jrvklDv7D2+YG+M2snDDaGs66mqjfrUF9BFCyoQP2F8g6Ew3TTuMJBLTxF48
JuS2og2qAswdPIp92ycd/YN8whYGienFKpYNJcuBO/xBkrwu1SeAUsn+ZrkBRvEZ3XNit8LIqmjF
mUps6F14Mz7ma1xhyXvLbgBWaNoiHHrGNHKaJmx6Rc9Fe7awO6ofkCEWyC0ijkLjgzuGH5DNlqvU
rF59AnQvrG7tK83F+LNpRHFT4GL8YVmv7ZjVunxwjYVcd/F9n9HJj47lMeHyP57xO/GHrV7XXPOQ
CHE4OUHyLCeVb1rRdajwE1ENst3eRqo4VFmj3FnGPaumBeI/rlPUh+AbS+GZpabj8hzrkzcFXj96
S80KRLvga7ENfh1fUolRlGS+1ZXs6ucHnbKFO0lfxqlM/5+zssq2LaGXFUGslf/Lowb2pXv9Nu1/
4TT7VZ3cEFBkYjXZ5C+qpHYcGR6us3PjZo22bBpVB0aVQUOt4SvXNVVarejz1mb8YNIjpqas0eIm
CRCrNh2VyY9C5PoAPXeIUTT4JX8YbmKJ2+UU29kdoo78DiqYyQ6ikw2oGNk/c673lMupqXAVamd0
6hEc0u5PRIGBl+dQgPouCAieUAjrgybvXtZOK+/mrUPgD167rIYg+uPkxKspGn/yENlhrvxoCyfn
3jMtNXrBn/yuYi+DW3ocStdLO5sMxzaW4Nu3JRSbyCE+W6se8lj/eQtU69kkHiJQqBJcc8g9Gn/2
6EL6wWAWYGj+Fw9koAEmunwjqs+03RZTBTPLU+FGoEner/Le56Ub9F+/6sPRvtHilnGNokMZxR8i
0qCVRnHsJ8GvKc+amJ8Nd7oKAsLy6ef9WMkLvlxN8/3n3WFgTtAsfiuOBoiHnaOIh3fS39S+Tm71
PlslisFw5SjVLvZPRknZsa+51QTa+SWArjZZAFUjpIf9mqSTmcqbPfv0/7T6uSOjqUO7+2mYbkC6
11GhrvuNTHK8LXT6YnYIVePAswJmXMZzmtVuL6RrEQWKrkDdJonSmGEelAfv8XwjsqNrwtyewHTe
39glbFazbTjib6YdsaOspJ3iny5CjV7/jQ1WW2us7Xt7hMS3vYxlIEP3/+NsaU0+eX3BdF97DWpU
5vScu7ng4/XE+0cTyixu7JzOm7lJg9KQWH1mGqgvFWf60unLJekQ46A1NF5B3ssyMJnvZGup6jHJ
8TLieAFiwpAiF3Lra8T6U6sFmGe02M0Ik2RzTcJAbOtGixIzROqwcE0vUjr5rqz5GRGwD5snX40W
vm9gqh77MXNNxY52uWItW0N/Af9l9XyEQGOrFIBWBJb+fL5TzlZoob74+/ZbGhNQBkKfoI+yZEG7
+iMyutm3vkm863ACyMFQXhyshdKRBheMlVesSbdnAE0IyEj5cgzb7ECSL4egTHo0QFItajexRf/8
J1TckKAaZQQrL5mMhD6uXkGvzP+RkMxoYFkRTK4xO/jIq9RdaXHwhBebe3b9xqC5+0P9beQpkYDh
Hr07ub635oLdPkjgZn6k3qA9INHVbVRhBlpQqqphlOP5Ir+WlyKbDXzpxFlEWXRiNGXRkBvVdzGZ
B3BqtqYLBWKpEpGTzTWqoH1wiFRtis2qdnxIGZXxt6Qb7jrD46mdlx/RC/ao4UXCNvgUYtw7VbYW
CwQV6CREiXredFMNJi42lU2fGI3+qCyrjEjRxdqksgRlt7K1+4wYOqSnZ4JtYedbDjNMrQecEd19
XfqDjSYOEPeevaDgxyY4VapCq+qgai1xPxtR1oyMj1Y9oEbdCS4E/FRKHEkPHm5sat8YVatqZYKF
8l8oPR5YkFMX5oX62+lI6vWOX6pnf3erNn81ns1o9HATeypzH5lUt5vGb0+VG6Hy5N+HIkumMosE
VDEsSpDsRdjfnnLwayFITZN7KBw6btTB4IH9thuk8y+z52wkTBcvS9V7Vd4WPCo9bpi63Qs4qfIU
79nwHTOGfU+/KkwgpdtPLTif+R8wPzg85u+vPVzdKvWT1ZadJoxj+dwbdHUHdyOSYoQDJk8Bohj8
BHQKLyXvyAx/6TZn2av73/Wy6tnGh9W3TKmNgkcV93uRl4a68Vp3TqzkflCqoMacrWD8DWEsf/8s
Ijkgr8f7v8SCqs5biF22V/RcSi1J+kOu/QPhXrdb+Pw6O+kn5RYv6I5iEgpU6dDzdmZa0GQkCtAb
4G9rdWUDmKUF7UNBhp3/bt9KoqR4OiBwvArah9r4EWzHiq1Ikm7jMtPMoa/iF1ECHxEsuJwa+LND
8GCru1M5Ww8JJXKTeyaXH/S8LAa+eUYa6ikOjeynpPy9sexJFWVnh15TofKKnapiQL1LfzpfzNwT
DBUWjFhbP3fpgzo6CarQ88q1jk2aRXVLb+wxI5POJ8UbEwfsl1ccdKZR0jg/HBZgni79/INn0H5S
D+gvmGnNGkRY0kXNbJwWV992rI7kJx0Pf+n9PDT3hYPzuP3Wcv8n4KP+DVKYXIrYs4PN0dptkG2K
bRNV5VWZ7rjEgiZKOCSep61RNqzBprRDndcJgUhUeSEWBlNqq8ekJDaNVc4k/ioXuLlZhsS33wGD
YPc2iTQxc8S73gJIFgBMb4CxtDRBCLhysDTXi2hHsSoUn0yIIzj6meg87Npgvp7viHdtovzjwqd7
o4RrUpp67PFr79YGfOAgtAF+xVka7WjdSJP2GSbkA2MSIi0CkEDYqRYlZNAiQK5cAZLSWelgqJHK
FSq/PwtRwNvHDzVYuOEsMQWYN6SsR60qZp1P5LbXiuofa0NbOCikmNVHuwb1QL0+tLHm361xBsg6
TKIf4rgAmuw0uTZB/OrRSYlhN9NedK3uP8tKYoQykoz+s7UKgjJrBe/oJ7GXtSL2IWKEyH2UDwsP
Hs+cCe7NDQN2q9a9IZv4lfaS0Zo4KzXlaeQTYyFmTiQZcuJxiQXkcfQpGl97giM5a6CooRg1njZ/
KqRrS1pYxOtqnWtiF/fpHG6M5xfBGwHF/SEZfstTtS9Oz1XDf4eSgTX1o65LsVY21vggyYV9ExBb
zG3xfgthNz/TLHz1qqiNgOJ3N87bx2BB4CuTGVlO6ke3GsfT/PcoA3uDZ44AhaHvWQxhbwcQxkzt
uXlqTno5PausSQODGT0u1vw3RZBHpQJTUsj6IeX/ni9t97vHJ1WB1p7KxQDwpViONjJWsMxUc8X0
h6+c31SYgcrTL7N3hdXfb8BxSkQHokKA7+91pQGNfI4JK84F2nKbqSos1p4NeP1kxcZv1CmTWavF
7zc/4PQUMdEkhWAeUJuG2pUyleB67+dNNr9ehQR/5V+yBIKw7S0KDAmAmS6EYZxjGvw/OUG3Wzpr
OilLS+p7I3K1xCgDAZv36osToFL4URFMxB4zslsx7VW3H4Ft62vvHHzqyWKSBm5Yo0iRnnUbqZDG
BK593lT5rzNQnzwgCv2aFfd3qED8VyzjWGtZFNwXzJr8lK0uahAUaJCKoUkRZn96OsC96CFxcHd9
4H/6RsLoRQctfkqrqeWc8jdcgTLGOZL7RQcajWkoj3PtPLGyHVjZiZOk55/lLKPCqgK2nCqxXneC
MvUKYA6qsrQ4VW/SzNAEnGw7SytS8em/dVlnJKmXQjGV8Sgt1xL+QD41++3VsZ1qylW9oCOYkqL0
tOtmQ+aMvXQgFCKd30RtNd+Y5sBGOJAEMWAnlJotEfZ275e0fpwSsuRSeuB88jGY/pq4vYqxWwoX
x+aeJIXNm6KbdfO6HnqyBkrsQKx14ET4iaxZOPRN9xPzV1K4zQ1KmOY1Li6HYbGqOq8SClZCONIj
fvqNdm/Z7f0doMxUt9bF+qrJtn7qSF4aLk657lCIREAIyAA+HMmCsDhUZLzRngksz20R7vlgxfGx
fcMMJ9/eLbm0YM2GaUYhpV4k3Mzz1qC1NjQBZFVK4OPt75M3uTUcBFlr1moIRvg1JPrX34WRHbCP
KNvLFAB+nIJx1rTryng46z8URCTyDYLqRNce+dZjClME7AsUMDUWO4IMZw8ooObp7Sr77YGT8d1R
4ygdqfpEM20T6ZMjUarLiiG8ksqbZja+fLxab1YHPaIiC21Pf6eIgrknmySUrj3CoGRQc7zd68Um
E/q+SSNfhLYIS/mQMlvmJKuLQD6sZOIpl/lMN73LzROtp77M6vdr0twG2NgtXSn1OynNbz8AEdWW
pOWQvP1PkIS9CxNN0VEnVKSFSL+rchjl/isH7WB8QjnM6YbYFpHD/QI/1d35fKch7kZLUHY4uKJ1
piVi7l/ZnuzbEKikuGyacSj2hAg9+BERFfDmTJlLdbKiPvzd1lE2qDj5bwApU/dTHseNXZbotPjf
e8BKTaU8WRcPnX+eyxjnY5DmUCWebudDlBk9fNJYkqeM6zL4DZ7rKhApaKUdMYILNIqum+OpoxpU
d5VoBEqlDrMScfFZ9LsXieVCMBDu0/B46xjaq913qvO4/wXmGIIoKe9ALQD+0A08JqeYZsllloIP
H4zx0YBD0Jx6B5Aq/WWcJ5IjgIn3hbK3FOtUI/DKbCoGQdBjLcPLq3MWFGDziJBKzbiwppnNTlGi
dOksTJn9ZSZiFwhI9KokKZ5mQT2zvfPddm3jb10k6uj5hqvB0QB230HsNZ6nqUwdU6HsnHSgu+FX
DLl9yPtaVZfVNI3ycJR4s3IEauFJB31mMQ7hlKys7LQsSDoIcBmTutCBk8Pyb8Ex/EK1xK6Rj0ry
KJA0MRmI5F8d2A0+uxTzcZRpvQby6l8v7Kvd+vnyUn4vlEo93UUOdMNC7Hx59og3YlLfWNk6+2ft
y3/UeXhHrm6GpnzwNGdR2UrkgbCXQR75Jn0qJKm79J7ZRSkJJSfDUtKa1IWnP35cu9gZOfT99AWG
nCHSv54AzFOLrqruc8IQMxeyLZJLEHzouryHIdmxVI4AjAHEfe3k7ewRemITCLxXoJt7iaQ7cPFB
xYiuKJWrKMzRNufUqTRferDnOfJ0hoFaDN4YYxoSlpn3M6Ia524/3uNMxgpYOeSbp/SMukFDe1cQ
Wry3RyKjLdq1Fvj1adSj1gIeMietbfiB3/76Q9zT/lGpM4tF3wTFjkDaT/p7Mq8xdK0semSfSsSg
oBoBhJwE3toh14KekVT/oZX5Qek8z3SMFT7gMhr4C6JV7IZkLRB0yhWG1L/7JLc5oW5vCS/YjITK
/nb2cerlgdbT9AIexgwXOqRF07F2l7aNq44Y/guzvX4o1IUCEA49MPECyaK2SCUHuGr/3KTCAnwl
dnkETnA6Me/UdkapbH4+TBLqBB0clzCsX0pfJgILFiAzs2Pt0724UOZ/HricasTdw+LfdfnGBitC
qIQGAMl4zT2EDivaBa31dJ3Ohox0MIlIxyPM+GfwrEpfbF6rhQGzMnQxDXXaVEhPm2ona49zPrYz
FjqVBWiZ+JOFcljbMl6APi/ASiqgo1aOCFDOag3/t9ReAdCOJ03v3yca9fLS78OAEqAZkkqqcUDP
m/GS82o8FPUqf520MaVeZ4fHRs1aJesD0F1lX0LRofatDyJu0bGTAcyX1OOVwkyCyBqipBD52vSQ
o/Sx+tFApGZqyMRcI0ohdrWWtqYHF/rli4rMG6rBBMNFmoFDzf/A9lnTKhNN1U4JoQGy444P9CXx
cAJLHruH56oYuFTeBl87giGK8B0c+hjVLSwSsst0wdZUO9sf1+uOgAeHSoM8G4x615yfj81KRcYY
xqPD6+UrHhcM0GLo1IbL5c5Hf+8rpkl1NnODBuDKh9kFEqnuRifONrV2Xpq3hrmXHAp4wUI3vs9Y
eP/0V5SMNVfvSnXob6eUczz1b3+Fhcc2Ycb9BkHH9nb1uGaDvvGg+5pgIApgpeUaEiUzbT/dmC6N
hI4mZXtZ9FF58LWqK4Xz1bjbaAI+DB5voAlOstiZ/Ijsqma1imnmpu4Vrzk9jSfKFmTXrfOiYq9P
tt5BJGcxgqowMIfRYWN626C38JAfV09W3tpL021PsWTd7qgqpYG8wLvUqfmKYfoIGqi+rk2z8Jm3
4taaWtWJAK7oLFWbpSK7B7cnYPyUi783hQsWTc0C4AXzs2XExNh+0lIYMKzi+Md/KY7BTRLsJn3A
h8RRmrf00WSFkKiGrnWF4beUdHEMQchjzbbvs1uGoFAqHIZnS2NXeiT1tblBZIOcokkzUYjGgF2R
mspwamEzqwOWKQ7/IVvz4eob0AIgC84ib1YEp7AVNCnxHg2JZCVl7nFjPChX7g5Yu2gJ+nHMNaQm
J4jHQT2giCcXOR4nEwjaquYj3ItPY9UtIyeGAxXUJC9L6vvEurhVr0k6xMrJ9lCQPoSdG4QH7AJD
Q//OlUENCVHhMJqVQuWlf7jDGi0o1QrVK69D/zQ2CJ3twCJeVpWSP2r1Vbjm/zvpY/pcsB40BEth
kBiyjNy8M2lz5SSytxfu7HsPkN2P+VvUmi/Idjh7ZfebtXpvCKH7rED/drlVy5q1o37kQWDz3D/n
gL7VSyReSYOHWacGZz4wwXWt8xEByhJdbYJhk3B/AhWM6AOm6C+k61buLnpD6Bdk4oSujTHoi10d
tw77kaHev58UhUl3VUNw4zO3NZZo2DxhTkql35RHQrnil+6ThZNyhRJybYphdfN8Q1zfMlIEiwl1
7/mvArVdRIQljwpWdA6ug9PAbgiDDdvxGm/v4C9GJMfn5v8z+dx4iS1vWSiCHcR+DdiP3OQN2O+D
SAEflG1tM4n6KBYepib/zLK3sc+MyNxcemHulchfrg8xamMVmZ0egwPfRcxzSPZFgG/FoSXT86Bg
Mbm0dn5sOMOiYcoCbXaUSKyaOC5YAhzweMbsS1o651J1aM2HrTi47DxTKSrkGv9WsHPyx0PzE+yV
6SUQ7RLYTZoNtwDUw/57PEYExFKT9p9fxOeRoImIroOr4OCBq6eTFdlEvO1Ln17dsOOmAHzW9uIH
WULl4yiuCj4ZskoK6IxxzNjAZs2KqJeQBGfFUH4+2VCe2nLcrU0uBFMgp6YnEVhLHoRZr/1C/bQc
1Qc276hpNo1DAXf+9AHWjb1qEI1LBMtG9DrYsX4nK7GEiGkx4UhC7TDR1HuY12kDW5M81OY4D4a5
PczuoNmxi4gvpghU4g1Dkaxyot5hhqPb6/QL5TUeS6+6Goq3fm6Pa4fVhNwXIQY+NEX81R2AofsA
fX1qY1ly63Bw0ksNfetKlrXtFVUOeqy+thLUKNALdT74n9FhipWAFKwDyIYbGEcu/oVugIivesCd
TZRzdsBS40mU8bnQUsKuBW7oKDhA2/xJD9SQz8tKEO2WtxLo5g+IzptYhwXe2HWaMkl4ExrErmir
j9Ri13MK0uUrv3ifsKtHf2sjlCEB4Xl7i8Pjsrg6SawiVmwMbDG2kzNw4ltuv6ry1vBqkIy/xit8
EJT/ZgRtUs4EG8Y/zKG7mYObIRurQLEPofff+3gVXe6mtrekGYha2PZEYyeCpFskhN6lACn+m/Au
geS614EO47JVhvT6H2ZoXXj1v6bAyCmiP3WfZ+DyHlwrl4Y77qQCSVXba+1EFW2iqMXSXHtFn/7X
ydW2me8OJgfEHsmSAc8K0eH5bYw6VemfKBWWI0C+KKoOyOxypk37RzMJd5GZte5fuUlBlk+IJu9J
TNLIAdWFp6eoZLY6phDJcxbT4YmXHSR7lFncZp8zApEtdoSeeGnWLeQ2DqvRFZk1/Wjzlhs5suJo
leiRTu+u0mjzLosnyrnCjvdvQ5ovvjTbIwr2vlWM/NgrjLFrgzwiwbhBSpD+203wDV2J9bqzThnq
/RxhvaFfzEV/YUf3LqNBdLB1c6f/TdrpTDU7fo4EOSsb1hW8urpM3xTr0JJu/cif/Ry0aDpofc1B
zBBxAqcOdXtV0LomeuDax09PNzQH0DKYRka2l6d37iyUF0z6ReVTu8RCZIOqY6PXnEJHtQwZc/w+
e1U7MRQr9KKL0W8GxZF1bVz7FPw6xVyaqgyrn25m8R7xZn9x8KUhC31vGiPIDY+6jNj4s3oqVsrA
MGvd+VWlC4EJDovSkqaQZIeBsY+K2ZfTgfsrBkqdd8GM5huKVDTDJY2N2ne6kLGM3kQp53zv934O
xgpqJgaTQtuGsSNOEy4Q27AfsNp+cP16FIwmg4R4yQYjVSG2KicoCmOkTnhhulgqRBzBac9Oexcg
1W4chhc2Q4r6Y4FWvvxvuE/twySygu/mkNJBVjU6oMtSuZ0z6sEFZTrBBZWxJuu0q3W2aB0eef64
mPGZloHdK3S6qbvOBLrVVbmtB8rvQxPxk88H7XE7MB3hQk6ibl/CrvAiirrBx3q7UrikI0hD8ew0
nduJhlUDUmMtNegBECHZn6EnBSJh7fZRMKfcswMNXO4JVUSbJsIubD2vKE0Nc91WaBEIsYJl3yel
7NNIx0dDNpLkrctZsumQ2O1+ZE71kZcPb1CP8wibTuyB0BswhmtV4asuz1vtzrH/W8Nn3Yk/VqLa
eTjMfloDNGib46EjQaNU59prgm8WKgouzTwhtyzX9Pfb893Pa77cl/mlFKFUKr8ajBhLblaqMIU5
8AVd629wz/DK8dKoFmxrR5LBoQysndELEsA+tl7L2fuWxVVTUKgC+KV+q4U5/xzl2t2UxssGXYrj
Y+nQwiMPRidHQ1vcqsAygOaTefwnUsRna8kNKQjt7kGsbM9BbHqeZkfo45xlOlupSM6XxJ3pHfIK
umCV5ieUmFcFK5oNn9Ahk0C7LjGDczXpMHAbjIH38f0IrvNkOAK3nazI9aJvR9Zut67dFV5oCz/2
8zQRxq/B46WG6aDhCFj4jCeLy/8jtNV02nodU1fLNIE4oCGEiq/88SteJm8+F8Aii9dWElSU/A3A
e2NcFhuw75G0EtYO0CO9o1BWo0QEedhU5bSxiV+JyluIM0G7eK6Pl0FFvBDvZChDXPo3QqDpSv9X
AGNfJ3HVyTWqnZ0YinChLsHXzKvl9YoJUIOJ1G9gFZHETvqcmyxzt+iivqh6uyc4Uwtl/Kl3teZO
PxH6UdsKICAvgjeZpoIA7tlNI05OyJRIZaQYTgXlNaWn177X5EBqE9uYjYJO8glfsnc421oPOgq7
kuhlzjche/O/98cn+VDcdv9EoGQPcJLOgTYLXCGY7abvTmDTr4gsSvFUEIeI9D60E//CmBVTK6d6
I7ymkHlfznlTj4IJvHRXOLo1T8fZX5/h7IQq0GXm8yluNH/1/SQ1r0xuQ9zgCVYlDREvvjGUMzZj
wD0CECTLOn3hjGUkkQuh5Z3y9mYURrlEw86Bu9xzEFTvz5BDnI8ePToGgY4icCvcADAb2PjoRCPz
DWUKxd5Ws5sxoWJ/nvTvdLQznKOzaJjak24GTsyy+n/jVRpKlWDUrns5AwXL3xFyEIeHaaXd3fZr
ayoDhu1zMaD66CqIDqsBWK06DwKK823zjQzJNLrYkTz8C1/OWqgvPAtHBd0QalZz0moC8YowfYmv
N89nIlIVW806m8ma/PXcCnz+4C78+gl2RVHOxvTlpRFsmCbqrywd0O0pNvQpUKaxfZgGqcyygvna
wAuI9mefg6LXEMV3Vw5WBw+qZYHVjDAHMWBt1oMXHZys1IP/YR+xg2p23N01guEXFgt22Ol/uVQF
skvBaj7X3kcR3SYCO2qiMgdhTKkZpzFyp9IxxVIKCqb0mwXUN3LJ2uA0Xs9ekfKE1Z17Y1Tu1/za
kiQc7E2PY7E4a6RARvYcNoL5ol8WxGeMr8zY/pqqmgcve0Q5g2omXPIFCgxQ+eN+3Ouwj2Nf/GNJ
dWubpuxNiXANiXHsLU1COmIIi99XVYseNUqnas9qMMrTCAB8cuQRvY+WNUguYkk2gvGIZsQ5CsSY
pDeTw0cJi1u9Il24gVIQYx4weBpNaegYAsiDqwGB7hXkljoUzGAW3Y29Mbyf8pDv3rL1bjCxYAyP
ABNNpFFBmYkQ4mpCibGWAqGaMRxBYgydKfAXF7MPAecPQkZL1pOa5wt8WAPkTwSGhYB3I+WJu94C
g83TkFW6uoTCPaoU/1iFgGm1C+ljxtk1ddDdlEzJB/x5bPGfZbaDy2OBl8HQeqdzVX7ADofr9LJS
mg96/jCeAAK0dgEcyGYrL411gUewvsj+PvyP5ty1PmGe6BDoPVVAIXbrvr/f2ktPGHpE7b4GU2Hr
C34vyDSCBJigwMapKNI30RWZy7DAi1+nIYnsdAaq+UDRc0S2YR38WdaAahL+6N+rSdHUWqNDqLp7
7Aubsd5EJkzQAzO4Pt+weJhwC1FqvGY0lcl+qJIrNrFCY1WS/yIuyQQJcWpEB6xhBHlGYRQzHix2
/4J198oCch/yaa50zHeUKxBYt6A1IQFZRyOWdNqkSV979LrEdc2kHAh6NEK0S3d17FF150OGYgbp
dE5D4hbYmcPxoLeSyo/VwX8Q3tnO55urZpoBbgq3bUrScXt6Xs6Bkm2JbVx8n1zUxmuqWTBE0Oan
daQF1Fvmu3q0i+d5ODphN+SWLCdat/dJXu/zebMwNmCkxk/bmP3Sozk9VS4UFqOfIY1qrbEZJij0
CJAJOMmLiZxPkQb/W3kVFlI/rd6BHqLP/93toL0jSYyRsnVjZ6YOpmTAp1PWUIBrJYSYcvcsnGR/
Jk4Uw1wRIrgQgfvDlmBS+3RWtMzmWjzZxQeLWXxpDC6PjBQg4qE7q217Wk/sEmQ8pyTDatteM2E+
3wwC8b8cLehfKQcuYAX/QVShjDe72ws1aMf6cR8rg7nIBBGRnoMQQnHwXNaZZITaqk2Y++T0st7l
V825tDCsoWJ7ymkqljagjHX12LpDkP14xsPiGE3P8T81PWfUCoFoQkejAaRSHPeYgMdlVxrq054Z
dVJnqJ45xRiwflZNQnkIvov5or/k5S+vWJSICbDaMz7Qgp/+ecYB/a5uvIOK2bm/Cy8MGjuPz4VM
BrB5rmmELYIFJRu2qHQhhTGTX0I6AGgxdTszVH5zAbIUWq//NzF20EwwIhh6cXc6e/gL0IQkOBbv
RY4BwhLiZAnHX/LJUkGs2ZkJn9atOO3QyBWknhU+7QtQ8wibkjmRJOoEjZm2MOwwMvoVVNBylXR4
xMffZ7RBLgxZIZxBVMFSRoVBD1TGplRooDmI7Uh1ZTUxGyKNZemng93Yu2jv2AG/aPRJThtNr8eO
HYdURPaLD+AFYASvaTd4vRugZVJQ0bf0uBaoFXPc+snC/HaQCSPw18B/oIX/xWopczVToy/F8Yf2
m3hcQXpnsk4F5sYV9mgkNbp2Xh11GyYgBqMNZg7LmSqWcajUhtA5RTGVhSoWOckBwtCaHhlGdHnR
mF6TrWv3EN3Mr79wFtyjmBsXpYyvpkLUbWrt89SQw1YRwZ42Rq8f4NAiZ8RC1WU0yGYek3ZHrMet
Mx7jZcq+4rnkq7di3Lfz38CQddjjvnNg3y8LtnJGTLKSTeKyusUDsFe9JGnUxIQP4rc4DtUh/lQU
VFb/nc+YeVAjCXkN0oINRy71xnFjWCIQrrAkPYPVhl2oKJmFf+vLOq30A4US2DBUNJCsqbEMRt2t
/c8fVbVDguaefze1waBJomwEG2qrA58/v+dfPDInHixeKUU8WQjGWei8JU1Q7Uf4LDV5j2qARWFm
ql4+whyuUsmFfSq/EFRJPQLdkXipxY4xaPKnVCLJAbj8cBdIcJPU7BfiDgIreGflUzcpiglXcwxZ
K51n2PvlW15orQiymZJ2z/cXov9XlrYJ9s5nA/PRw7B/URxjl+qudYGqVM8w2wRdLMCLaxdPt8Gg
C1DC7aEm3X3/kdB7NEKYPn9BODI8t3k17gUg1D3fqIi0TlABbtay00E6I+ptY+sP16zG+IEbhHFo
HHO/7GKx+onzJcYrE9w6TyS1nt2PGKAMpMs4YKuUu9+wQWd703r4ByWRpM0voRsdBx7rl9efgiDt
XuHWMU+cr4EDzziHrPa7zPqgFoDgBrm1rkTyoYzBqP8zMN6x9R55XE1UPA5IVpHfwg4WzJEwfq9r
K/wmePn4HOx3iK6vKT99ZE9R/PV5GsMafa/NbZ/phiEklccEnA71JinQSGlHjC3B9xCn7+kH9YKs
47DP3GADZu9DD0RdCvMMCT9GxSrZC3GhFaMWOgI8CcZnO14ndTlUwAKNQ8arI/JdEfHZTQZKDFXU
qm58wi7IsTQKjb+k9sPaa8ZzMLMMviQJx23rSeEAStTg+WuxCFo+XSDefWIXhDizlmUm3Zrozd+V
E4p7o5o0bH0mKl4WGRrhwGu+H+/y6OBNNXlu88Km92z6PL0sBxfJaKB+dKmIqC4KVcjXn6Uh9D3I
50YcK7Bpe+0+Wg1SbfkDy6Dd9MuTwM0j4mQo7Uwazg5GtivRRP/2AXYB7EVPSvUUd/PLUDAkIfa6
BJgrwxkpiWpPUm9pv/hJDaFkLigFv7ZC5xqpdgG8ONiYOKS4SEx6h8Cv4bp9OEzQQDVTPJe5qtbR
TqkqamYquyQ22z3zRCK4Fm2joCX6ecEzmmlfSDwtzYcUXBaDLDSgsc1on9LPcpLQeqHipUWGeidm
M0oXtB9emP1SGwhRfSKhev36VWd8pON1pX8K5YmOtvtNptdvsvNLmqYn8Fj+w3dtGF6qUybiDsoa
Ef1UwwMFGTyln4HQW7+wRszpD3g+EbIzo/+I16AgG8kh2y9HhUUxab9SmzjwVu9kL9zYq6SWvR9Q
uGVulcPhAQvHpOnTXIGAjdCxEax2ZBic2CLaON1BjFSxli+wXPOS7bNQSLqDGbL42GVneAYg4hBi
MWHekVML/3Y0BEtqV2J0Hadoq8Z4Dk5bnrgDpHICIQHJtumcCi/sVgVgcgTNZK8jMn8d9VWcij6A
uxnpN5JIEZcCser/jRulck7Ws6ehzTcimbUm0HuKVVFnHnNUavuXhqlmHvpeUo0lZmGOZVPSfEfj
SO2/vLkDvN4xb/6fiINL/xuPWDXeUjSmYfDG9ncRO5NCHp8nfbdhqaUDSYxCm8kwyukdmc9n00Ul
LUTr/Y8qeEBtw0M1+/aogTzsWTk6biNYjAnHJHwq4NffqtRIiTd/jmbCIUW87kXj4un48tVEkDNo
g3Q+1zvlazlLt3YAIckm2vojtw4EdkuEZF++jdT1/8IPjCdtCN/5S8Mefa5FqKRdhu/F2aOyvWmK
+bM0gOUtMgf8S8hhU4cOu7d+u6OnoBZtJ1B2L6kw7hfUINkkpUTdx2bA1wL9AYPFQ7Fs/XkPe9OM
n6Vk5IPQm/rC789nnWc2bqprj4a2cRIwggmxB0I8XHLL3j4lVHsqyb2UgJjcdjjOggppnPr7kXo4
FwwoyjY2ISAl7yqPmsJHJCC0Vtr7pr3aN87qTE8l872gRVxhGMKRVFyn+VCnMv0HdOLeYgqxuNVq
vRzD41EBTB42tEDmbxj/VDY8OAB395BnuyoODhRHq9go68jwJZOZPi9IZlsKbyJRsIo62wFa4uzF
rqhT7eY5QZ6nSBMLFKoIM0iNlRhlljgtlYh5SKijOBtfxMo/UTm/5P6pDm9rj6mEFFdopGRCwDVq
WzmonedZ/CpFp16MYfsNLSYCAoT30keSsbkqgocG+dHr4608j37aqyniT7k90wMiBPBG9Ka9g1K+
lxpibT/QC9AXJ3i3xQtc1GZ4WzjmOrRBiE06xgLs5qL3JmdEUIz1oAMFJcpbGs9eS45Zz+tD1lK8
7KyIiSF0UwO/AY14GZD8HNxhtJAyK2RQUY3wC9fIYpV+oN9Qw88fgr0uoCfGxKVKB55fmVxxP3Ch
Af9CErQsHBqvDAZLPc4BZItAd6lb0uAMmmJ4IX8RAV6Oq9leyzjE58WlybtonCt9BjOEvQy6L/ol
4sqOEztPXwYq7OxcH6rcvqKzKQqn9o72eAJzBlQhsOlXBH6plcK+VKOd5/AWSvJrWhC0OHZVTvmq
Zd4vdYq8yzEZPAHoxoNc+7W1jAlfizr+9KbRcyfFNbx6CjLybYR/1kHWnb2PAVouKuzxRi1Bal9U
AKm0f+DBeVHH3Wpp6g8tPR2XzIWGUE05JJaGJyS/issTIf7Y9/+55ArjNNPu23lkQN2bFBRAxn32
4Oz5qXY0aBkpt2KGtVyQ5O9jjskeKNZLWV4JzDQxQs3sQy8O6jpQ3udv23LsketNFoIhkylVHZ+0
wny3lX8Ts/ZPoJw34leWmM8MwFkeYSeWP715S+SxL8n6471bXOFrikyCE8JZchJ3l4tk1HmWQJ3o
hlizN/hVU8HdLdoR2DfQ3YVqaoHwcJl9K8m7qk5kN7sVxexylMZJsaXTHBmnIqNLb6OtBPsmt6P0
oYsAMQhcxuJgkQRyZPTu/ZDEiBHSC8EmUNCty9cPjJdMnh5Me8z/M5JwBEVdeEHGnAss+kXxVd3a
wt/lT+7tYsgdveTT2bFrmSm5TT+AnqhxP8PP49vV8hKXhAFcC4ltrntu9Th8KRf5D0P3tOYxacaX
TA2vORkE5yKQqKNkVDOPuLiaHB8sYUjzZSLvkPQsQc8zBtyMYt3gfpXedc0HXgrN6wEsUDAqJovp
WQr8B7ufhZjo3Hj2emvEm9IY200OHHoCXT81xbVkHZsKQkx+AgM6BRT4fFU7UCe6H7jRaKBFJudr
5FVMs6hhQmxfQ8TvNYFPEYpe5TtaRN6hlHIjCfV8i6U3biLaehQjMDNLP+faEepGLpmhy7/JlxB6
V9xSR/aqBUB7AIWwGHs5UpxQDQ0mVOi0wmbRf6al6V1E3nbAgftnRrtNIIW1s4Y5po+qzNbClBe3
OAdoSfAk1mO82nQBVTw9tsVEdPJmDxxbOOubm40Y2yOZjUr/+zAdOqMAd0bkhQi2Yw04U97drghI
JCDcrofFxYTrb6KaqH5R7J6WWUdqAz9qJmpYxbNGdP5lv+EDJQXDHYFX87YhPbNINRIKOg/2x1Rn
3u3PaWOUU1tbXNwitMnluQvwx+r8KuAJv7XsbDj+n2BN6YenQUI19h4fbUXPqbPZa9RZotpnoukh
P7E0qsrx8c8u5N9le/7fP4xwDtuMRade4enWsfOQucXt6najV28xLBIK7ivANHnCcIjcFFeJVjOU
GCsHqgP5CL9N9pM556xdB8bdgrBbjR/U3yz/BPkoQGXO/fUbgvkQmnNUyjVDKFGz2EoyUh73AQS3
FHeGnYUrMh+McTIytkng5n++fQE87dWviZyrRO3kVJzJ9QVExj+rzABVtP4scKcins+8XSO482Wu
FhlObS5+AfemXd1fgnYcXcEdnrKE/RMGqIKP0rifosBb30DHpO23+IJbQxeX/ub3q4WlHOVP7gQI
TQyGII69nhLHj51xkViQU8c8wt+qpW2pygp9VurcuvWpKlWta4tBazepbTMHIRgxo0t5F4ISt6U5
KVz2lhn5ZkrXeNRJIhQ9TY1ZW+6a7kImMTw0HiWZeHG5+zmEVUQYeGom6fNcljOb/c2Ht4V1q3Jq
iWOizyyQw2YVYmHOgfIHuNG75bhcnElzoD92L9DqbRMPEzXKJBD3vf4dF84bgRYE8hflHAbwqkBa
NRVcwYgtKROunDRhzrDzOWPJvlITBOPT6fbizSWe/ep6a6+YA5Yz+Z69PhgztxWdLX1G6f596ysl
FbZ2ncTdfDhqJMFWe0ADsQQKESD9YN1s4R0fPt/dupx5CNgBcGmKbA0qpakK3nwLRlT3wlPkeMsU
Ej9410LGrXFt35Jhjg8hZex3uGTMCKbF+aHkG17uw1mhDqMwAD+rwlU0RxNNK7VIIPWW5APQSvFZ
OOgL/yQhofFUahS7ALZomcysI2sMpbnUwyrHFdp+vgo7YXAGt9C77LVyesrkC4O3l13SzRaQlvVx
x9hYnAdCJkwqfW6vCoTpDjZOBhAHlR05YdeHZ7Usi/p0CKPaooOiRoG7uihUFMZjKaluNQb7juWQ
BND8Tvodnk5cj7exM+xomTXXRTO7UIDEG2Zv3hnmfINmIqfQp4YEI+yIM/EfaE2bPRSJVZlc/udu
f2pGvxIejrjrJxujGvBB3jWc8AwU36ePCrdnMb1jP33x8jM4sBkUS02W2yksPGRi1wJE0w2HAuEs
KJkwVmSHV2sMgnOpGrTEoVaW/Oh32yvjvl9nNpMiva6fSoC5By3HLZEb5Fnqn2FgO2SyMkCdRQQL
ky+MAqsrvtsxItTkB/dWAudJhwu4516zzLdiWG54V9lB3Da2QY0COmDSCE5osuYxNmV8SuvBeqWM
hpv1gMSVae+Y0s6ksiKe4k0IFGSWR+zMA8wdPf/MqYWkGeZ1yW6gN4O9MrIyPL8fnVmiiMB0TeR6
u46APEshOdXVQr8eVzoiI9veKNtJFrbKFbaVEiqndGTXKJn4b9AJhhTadH3gjIfdqO7ulhYP6JYJ
ZdFSJ1cQDUbEwTKm48qTer8tbSZ4QjdWueShJY9dRxoAEuhPYdoxCFZoVTAnJillZDJYdyA8dyP9
9vV0agoG+bXfUbI2syR+ARYBkGz+P4FmR5Qo1tE06v/qcSA+fcJ3Ick4RmoEKo3+LZux09Zi3DXZ
DLNU5gjVsETOWK9jKttkIbVuyJw7AK14fFeg/jmiWkct6ucgwOHZv6t/5LwQ3lzjMz7WH+rycMw+
pi6W2Ky09rKZENaTwAgfm9Jn0B+/W6K1FajcoORcO2CeqLYjv1a7pd0Ajuw1Rh7aeisYwwgFLchn
4qLDvFnOLSzs8CWZcLPCXQHUDS2j6lQsfoJqYyWd0nKZgpzdMPBwZAuObRs4KfoJwDdOKQDBhlz6
33LbgoM0yBW8heu+V9W5OtxyG7dDlXzZ5sntGERVvaOTCMGB3Gqe6tXsxU7n1z5t67shCUOzIOAc
nzXi/xc9Ewt4DJP57LgucOplXC4VyALGizxVb4x1jKpM4r1Rk6cc/t1bxf7mGUTtwxRXwHMYHeTs
k2t34Ncr1RZS6Sbvkv9yS0mG2UmQc7vSPtEJrzKDz+zjECkAY43m+Gzqh9lE3B5RfGmL4eLTumTU
/5d1Ca2Oq3UeXBFm463BUsEejWBji/3AxmSkAIW58IM1J2WOvnnjarCu2NHJu4xMCN/e9zYctf5m
De1y0KTMRtIAKncjjvpDmzXnXWF+RMHUnJ0RE8yItMePIs7BqQ0amMX7D/C8iUbe8Y1cQyN5v40G
IeiklgRLwv6TnSpe9PiFI44ov/p+smtQx59ndKh/rDOhGSsgqTsA7k9iPkBaLpskBgExCquxRtGi
imWTUF20MtYQTHOUDkt44pjv7W1mixg49qE0rMv+N6B0SnMgUU5t6yt9A1d1r2rUE0JC3/Td33it
08XQ/EI88+xloer+W/oV4YAW/8gFV8arWUz4A1gPx68h1Miu5A6Dp+1o3Qh6JBRTYsJ+TMlTBSdZ
6aZy/FPizXMBuD8izy5sA3KbpntNsNjx4F2XRwz5un8H7/T4yewMB03qiDW56Z5zSYjm44ZDGiZQ
4K+fK7Bj24v6MkWMXc1+fR8gcKFlBISlv4/T8dOJitpT5PAZYTRDaAmAmz6bbcS76DxRNJwOai3N
hTIljAO3/tnxA6qVjs8BH9N+dCT5lb2gWMnCmJYMBSdMsIRz+VbEsdAupEjqyVSeb4G7tB/TVJXZ
Z6+tXYQlNruYM8XuDsLlVVfUXZxHrszmJGzN8Z4izyeMrsGxeEfDpRuesxeDFq3aJupeYhR+BHbX
31lB3B/Lh0dgIaTZaqg/B9V42VNbJ3zI4y/Cd+iEw8DB3RNwP0VSqqS+5aIgwTYxZtd9+xiF5+D5
BEFuNVBnS8g6ExpyhVmCID2IjPt3lUtQC5jOGvZDnTbg5ugA6WC1W0GxAOUYcfvTfp/tqN3zcbn5
B9X5GCc9CiZOyhQ+OpjYdW70gg+PtARG1jBevkOk1mWzkCXUiPDg1Iw859IqSB/hMhXLkLMG747x
7bdsbzn5MwjO6xLaZ6+I9/mhOPMDE6Z+QLgQLFm0c49MXDGN4PRDyXvCO7+PYkZFSMb2D6DtYi/e
vWjAnbqxl4qtQLXUCv3ftUPWqDrkpH3HC6+ZTI0RAVD84ff1VzXXemTbpG4W+9s2/lMMPpAIYyB6
6blnecTa9zx1JEo9m80t7askDN8qCsg6iiu1nEnYCTtkNMNBTL9z3y7q6AU7cFfCjkQKoKibm42T
qEPnRajN14WWUO94iULKQZymrnPg7LNxmHHa7WTkgO20DcRf05SChiEee5JPRpOvTk8Mg22AW67w
3QnQQlSfezdMlXChMANQ8GvOgbnTV+Jop9Adbl2f8g18JDH/e14PgeX9k0MESyEIxZ8NMKXYd3J9
8m7M5FM7v3Kffc5pqjbtuKijzoY+N2YvRRmpQX/Hc9eyVDWhtfiJwLbv/Nn95iNiITK20rE+NZxm
d0AN5/eLY5b3UzA+zlAL6C910/C5WT6xacWr41KNCG5cNqtWkW3xJePtd3O2Qwxy5Nv8lnkz4Zob
3+loLaDvvoNTvPVbOllBuBpymKgnInWNxNhyjv1HFIpHabJ/dfXsX93dwlETjMZhRiZWMJQkhaWd
iccr5r9aIfKtvZ9buDqZuFQeAW0y9vO3rnkuQbFAQP0ln9F3uUerMY/fa06mvVBw7RsCyXWcvZRX
ze8xc86xGJIZwYkY4FLs5jyWoXT2fXYatUofNnOutGc/y9Ay5EJhdnLbxmZcY/CC5fSa+J7+y+/V
KacQ3NGKMFY7r1Ymd0m/kwxonh2PFq9qOOkT4k5WCXxezDOjLtofPVIRTu8MlluMOAK77CBa8gUo
tAp0WF8ENYv3wmsLhuvPfle/bh+2TQysPiCjcuqMZhuxSEdf9KBXYFlKbr/gh0KWILw1x9wtYOu6
7W8NPhoGK+FJg8zDfUDuRowfq86orfChVg6ZVdEd8uLVuCVLTA2aKBygI2Wxyip6xVUu+ZDdKw+b
N8bCfsQ9w6SciVnlMc0VwF31HBCfoLh4i+MWzuuiexWlPdYi/02obO/j/sg9w3UGyHSbRpJqf/WD
llW3i98kdzRVKSP8c6wtbWWic1IUefjYEStUPfkRxG0b4+HY4gkKai040LVkTPhZnVLDE5y7M927
T3Oq29d8eh7LHD5dercEPhHSED1vborXM8gSPVzJ5vXOZLCam6nzTwpdJ4/u5RlY8ede/w9HrWF0
gfo9ZRbF7nvc8l9wiqjsQAtc/gW80UhAhWurj3KkLnYCc49awG6KmtQ06Vzhhe2yg6nMuPmWmamr
Lgl4vPf6lzt0zDaERwOstbJfI4tpouYixAz6OQ2ujKnNfi+kenwU8fChGhO3gld58pi/XKFp9uG/
6KjOXp4waY5gx1FPZmskbQkljHMuQrPAuWhKgmAy50WuVlV9FRTG5I7LBIvpeW1GV/ZjzHNo0/kQ
UMmoOZsF5EjHBB3dl8+vrELprte0wiO2+iOBIp3z5kr1AUOdwvpAUn3a81LgyvUOZbPH4aaKYX6Y
kVn8zwmfO662qMhtfWR37nKl/W+OArITAfhHt2tJi89FQhFnzlbb6iXsMyilQZvfn5iA59IJepbI
sHYhGD6HzD4Yd0eqnKLyCIIB64pDyiH6inzVaeyazOK2glF65yUavuJ+1HU4oCDif+oYOtaqQMJe
Dkc0DD7Rx1E1HlRiLl+89ez6yDLCs7SS66GFW34A8Hak91Wc6Av+cQ5V9ZsPPegAdegpcVj7L7Ig
GhB2L3PNKAVdCtRPC9U81GQWAiNdVbKJaw4oQ+ftYHAtIFldtI4AMoayPRFf607iu96AFWw/k6P1
790+ucyw3aB8KHzZNrnm+mK5KdFfdQsBMAhPnxgGTcqSJ2X7vLVYyvNyfEWVvjxPKuKlXBebTEVu
DwJd3sfpS3ung0NSVJ/3/j7HqIy1Q0xSaGk1pMEVsjY1TtbQd/B0xDkE7+pUJx47XFNBysutUWAQ
pv5y6XsaAgkGVTzyYDuKN3kc7ryDF6u5yNaA7X6e0mO5eAPHhEJvfZPVUGAOCpDMxlWJBqHecGmA
HUVeAxb7zQkWEpCbSOZx+NCMAsxf2Tq/WiXTH9Kggdz78/ImMOb8ozPOCMsa25cMtbn7hkHBTAzf
pYemFdXjxlZxaBsx9QaVOmrZhPA1Ps3NhP6Vl6TBdJsi8+bijzlBtgXKfJ0gHkZogbKNWbJpzqWG
EwyXVCVX8W5cUGoEpQhX/4XSc2uuuOgX46aC+H0PzCHPq0Lf8hgzDMjTwDo26XTNGFnpAVJPZ1t8
QCjTSrRMRTdDvtImQGAR1gOJ5bR4vnc2rJ/G0iCXDsi7I/upCD47KIh8v6e6wBh+YeJJ7i6x9geD
fDaXwfLSxN2bD3EHBSxAqaM/XB6L5ZTsYdAMoT3KsFpjuCvGbs4J7qGWEs2vmVLLxyPGsUWsQf7J
7T5xJ7QfdQfFvgMv9sD8vhO9kB7iBr1Kc6p7ILoDZaHHCJqNXWQ/Kjn6JlOzwaEgJ0d4kEEvIIIG
VhR8NnIjVQXQ9UnhkXVBkgRwCT64fadddUwaXnj5iLNu+RWcwomnMrCWCDhYZQr3953hT/zch2Cm
HyBTosPPqrVhFqhISe3/BjrZMjBw7W3OjqxHMC1Fye8V9/f5CYVFzCofxQwJEVfqh6ZdY0JWdMWm
s1jhz3Ck7CJ9fFtSo8lhejBHpI/SuQ+Dc3WyMjUVlNF2NjeOBd7b64WOwIjJugxCsGdcJMIVCH8o
+FSZhTBnBR3jmMFippJC9+pUkH48nU/YWSFUeTc8qLZobz8HS2TPQd0EX15pakcS0DG0k36ZONaq
v5Jr9CbCoBRMqZuDFwazQ1ddvMhQqgGcMIG9UuYBhy5x6ov0qJeDVABnazO2RTaYpVrJ6FXHrB0+
0QVxNhRIFEkhR+zCxLCbYY/X9yM1FtsCI+7n0QlXl02PFeEIj2LBsO2WwcoENJEUX4XQbHX77Ppx
lh8DqBwxaDjn6bEKthPJpmQCrsiRkLusxTQHV77NBTQxnbe5ZowlQVTCHDFhb2zsORxZWCredJ+v
VZdvp9GHjM4LEkwpNcnRx3PV8luvvSFeyNVgoaC9iQDPTP2fLN4OjwGy1Vnocmu2ZQnh+HrjzO1X
2bgc/aSSwBvO//1xu1ipBot0iKcLSJtlSBBdmdFr9A1Zu86c60BwVO7Cs/jiTlsGILXCpo20ZZ5f
A7w0Fw33CDsjEkA/TQthCidX0XF3L7QYboopRl1UgviQK0rSbM/jgNRsKfWNMsY0NowBpSyczfG2
5QbRBf83AMO/qNQI3fONCCK/l6VOJjxxR/+e/luetPgFbxHorWkopW5a1cJYcwYMgYtk7oow7N3a
c4YQi4051W7dDmUyEM9gKLqf8SwgUMcWinViqfNrjvy1G61v+IgBvZhvblgR4zrtenA+sAilz9tI
aHUFoQeA6ynbopw2F/ExggsxJGqa41l6VF3JjYPoOheHFUh1kw1RoiFnzRJOwuekG/HBVr32vZdT
WAvpEwJ+BYpna0bHLlmPTmxPIaAuaDaHYau4al2aL6KcaDJpulY/hk/TZWSHUjja5UMFRT1uIh6V
7kl399t0nYOu5puTFrv7TH5lTFeFQhrfL1ad1waPR1CTINEZGAi+WjmUfVoecIbCFvToVyRy51Y2
YyZXwSiPM91PCjNpc2rnwsuu1hQFZRROaa065KJiTQs/7LEyTjp3XaFy0i2HAvyoAXtRbMcRdXrp
FyUBUyF3vpIz0Nc7j2ckHj/HttBdRrzM7fkdZ4bCjC32vM52D/wJKUxG29UPBrPzPHyykcjhG7h6
DixvwCqHKEFvgj7adhydbaV216W7y8ciCLfuruE3DBN72UNHlV8eXKPIl+Bj+AvVQYsVADvjA/eT
HF5IH8mwA7UiXiLFXJR5RrACEjHTxVja5Na8K4sd+u1aQ1Bvpj3EcBB0wt6bLXuJxLhEiw9OG3K+
UrmpQvOBzERqIC2TYmGb2y2qyXf7b4Si44bF+gZISDpxPx9tSdEglMD/nPSdSTlXYnCfBZ+I50ik
u8QmXqRUp1dmaKveaNyR5CN86PQRMDTnd2E5ZwTRln+VceGdhsIHZglUL+nDctUO23IDluMMaqnJ
P7lzmmsZqiZafgBbGjLyEHUjjeZr/EhXLvDKOhRbX7PmF7wdiYgzttaTgW+Y/wOvh90JeV+Uqtk0
iSx5QLLOG49wkBzORdroR8ytKIkLmG107mCofO+YX4ESrUD2YuEKEiZou+ap8OaDoqKTEbkS9QTQ
hKqKx1SQWaDbaqVlqpdAhQN3wHQfUY9ZFt8JIR2X04CA7wud6SCZbjy8j1Q8DeOFtLZVpuN3Kn3+
r6zJlVegcBEXVOphg6Ne3aAZwB332px3frZL1dlnX7ilWo0pXhZ6lgT/fRPQOB+Q4uvSzr5UTHoK
gMEyjthUtt37LwWdgufl4FliJgqQgiGKaHTHQKteGQOLqaNL8OSQUkgfXDMPSgP2zHpfSv/H48uy
1QndE2EoDtozd5gAzXgvA2xgdaToYbYFQxPoIvhm0P4U9nf6iNID5gWEMIp6v+R03YNRj1AFmJld
yJ9sJPqI0sA3MrWDX3zhWK8thOtuAB/OvtjcuNhoEsYl4TjeZ9VZPxYm/jkQXe4e0XgDvyT4NCgy
0JGvgCT6L4KolywUl9Vy6stcDhIvO1p0/hIOLOGTfJVp8q93z/C6VIoPZ7lKRjweh0OiidEDreVf
KvV1RwG1uwXO/lWW1baw1FmLiZauoo8zOcfULISCpp6GKJ8IhmWaSujS+kXOjCM5UTk46E4V/EMY
x4kYZQlQE/iOVzGw/iL/SmEYeTvi4V8ERfp57M/KqtC0JKk53s58KBtwL/U9V+w1KsaI+8i14nVO
J+uDMW47UWyNidgXqEG8gPp0r5+4Z5egH2maeiKL+4KNwhKkvi+ebc9nlF0WU0npZN7PPhNElBv5
wSwBWyz29KIAEhXYK8gztLojnDR+IoXCTJjGwMsgLGyJG0EJDdk8/I+6frPKhf10W+igl0yC2DPu
XnE+8I1Z8C7C2ev07De2igKxTnw5QazRSAhXdA2NGiMlW8EU2NzuU9XUrR7srLn1MQUafGYJ0XW/
abLhArjpa7XzZ6XiLOsdGiuKwcFVMDT+OpOCfEHjrKSaq0k4TRw8w9yZ3gzj3MkHOOIrkcg7X8Xr
wnWFD/J7xa2lzlh2zUAIn6L4NJTbmF44dy/kbwY1fAcJxEiJTF2oLShs2tz+JWS1FxAnlIwM5T6h
nJi8Sp4pVDLn54scU9D64pj/pDITt5fRDdejdoLN3zJHsLucO/NFLw2Zse/Ij8xi0K5iRmbGnyuy
0dlItxNiVa7Hnyd7t0hxouT1rII4NOHGk+qzXLB7lMigNz1HN9TPJUTfckE7VMtYHjntO4M9bN4c
vWa3w6R9ADvZpQK5EWfheqlvRve2sV35kce5zUupWNLv9qbWWDAB0qu/peHXr/0fiGDjfL7ecjSa
j/5z5RkProQhjhvipM3ysojiaZRcaQqMRTEJDrdFuFxAEm2xLcH7Wtf+rzPw5Py+61RCzpN4537M
Sh9Q43HCu4TNTEulN5mFS1H5m7hpeBtdEElRvqvtwvXw2EpNaM1E8uS8Vjx+1ISGllxVYJHjSrmh
hwij+lDX2f98AXLRr6YSyhJFbVOJ3VfkUKLGdFjX5CKNL1+9UIrpOR18XSJS3Vg5nctKjY5ck8ey
stTEg3dunW3nVGmIIHiCiJ24CQUrg50Ov3NLoeO6G3PbeeXeb68HVti5DwLO7Rrjb09Fts9MYvWB
+Wi5Qbl/XLjguPzlnPZqyIKis/k2v6mzIDEf/bEJJGlGrYuHP6AqMZUrMsjnxXkbMvNllWE2ToLk
OPrvHj3Ncm+3DoJar9/Z5nSf6gENFWhpyRXBpdPMmiOIOuY1bBhSzOi7sM+uLkY4aA21AnrXB5kH
IdAtZaZch+ldN90a5Th2yWTKPx42yrt3ZMTu9qQx4f261J1+Dh/1dAYOfkSGuEVXPvLmJfobTCb2
iOgIbXltepgJz0ub00QgoSqK3fFz6wpMBP5S4elHmyBDvgL1je7mvt4GAvcqt3t6SZ8TJN8ybLZJ
M/mhcdaOOebINonHR3OwbyxXa5HFxIfTnIRpLajFDktDCHXh+9qSJOXYdy7A5dETY2DpTISRraR8
/CNnofodmTQULhqHQPA9yqk+7vMmKL9Wrdh/NPaZmkqYZKVXaQDDV552JNN9CoFiLxH6u6y/ugRy
oryxNks5ZiwMImPpuybq2kMtvi30MITC3UZbupOAOfZRque1jCbKavrvTZXzGlXcE3TvtHcXqL8j
x0t4tiGU+K7yafZERy1468rZN6L2auPOvzepe57c92jqTeuahKml2XCbn4n7JjfI2wHtIr8AK2r9
Cpk8B2jSfmrvSnMiGm9O4XeoiDNlm27gGgK9oOrWd+fSrFAsTlL7mrL9pBT0tmYsT/4LBTOUjsvz
GpIxEsyteXlQH79zx6BYz8ReglG+3zhKewm+iEqr8ECjNkNlDXGsOx7+xJi/5jIwgfY9gWzGxtDD
X5H1AJjvuJmNngQbN7sT1qed1jXCyTTiGJ0jtoUQy51aSzktdYZTbbJ5aYFGI3ytuktMKnm+EGDP
6k7ry9UNC8gZx7rhwXcS9fvqNkjyVQSxA05AaUMdMCDYj3aWXFDBnAdA0vJRu93P7osWoJorKsw0
WoxvX7AP+XXIRUWYYi1McEO3ghr9zcAPMPO6HRqhWjanzHBLFb61xnSWFhMrOwhbYdhieh/2gV0X
VDUbEh/tQ0s4t9NAlsDPh3wXSjZmop5SNoAcOuQXpfQGWPZJDoysAvisWPZICggscUFaqpw8Nn7C
mzd5uq5u6EXUzZez70Epp/WtJhfYBMwpWGNL7lBO5U4/MC3JGKI/BCaNTafHNARZD+ghq1tDeV4R
Mv+JYW0vDBMNOvtfjIMhQHn9kDUGSAH/tP4tEJNnwIZrQ2cv2It0+wodlntHZiynq6W/n5YBhmTO
Q7y9FjND6xyS4KAsG6oNfLtUj45RHkE0XQAelPaMnQ0Jpl6jPwcTru5Y6Vi9G+HfESuQ77ZBqplY
s+pAaggkkGt4wgMaGaADQexIcC9wv1kuek3Bddue9UXCUWTr3bioCQNb4iV/tOgVdnF13z4skAsL
jY3hwBsM1bKXUzNAswA7Nq4PDyGRUy6A8IeZrIg/+jzmgTnMcTqSamQ5nyue4zeMfLIY8fSUjFgq
cSvhkyeBihALU7FB5+i7U79ju/KvPFvSuq9LUBFEhSKDiR5MdLe5o/mdxWL13CbwP4R/8dXg1/zz
iTClevs75tL+E5L42qA74hwofaVfnxw2riw/K2MpzkuEfoxH4ZkRCtYHkwKQ5INEI8REN3jpnb+b
+ETBtDUwf7jG5VuACokfZ5jFXlM4f0YDQmzfC2sJCAHRzvNHMvr/mDqYZ9dLxdZXpfw6jMssQvXx
nq7/mAq7brqS7k4Qj4O7TQn7uDzA4jDx961iBlQ1ilrx+uYfZR+Kxiha1u7l9QaB1vijZJC3gOks
uKcDlAGlvsNF4tmeYLXgl7elKhqVIZaaH2y8hBhD/AYhzVkInlJ9S3VRwS2rrM7d713Ir9WXyAFn
4ysOBuB+nxXkFl/PQMOI21287m4ltC1fncP8dtcgpxpg9IIoMLgi9mkD/65ewmHosJXLAYVfYbbS
jP2nqMGG7iuoRuOYBcIG098bS9SBA1SVxnw7ISY9hTlZTI0f1oF289Adxx2gHXrPqFPhLe4eyhU1
xgMFBYij7jpZsXVxKUKKOfACFJ2NK2KLIrFOgmneOFs6gE5j+fiTgUMpnjr21IzU5dVRJY0N7KGK
k9VqtwoSfTfFS2H1XbgvxIo0FNX9qsycLwKAz49Lnar5ziBpvjlC7RbRJP+jh3Fj1RDpwdjXYnA6
FP8lY4uRLoYGoYOwC5x03v+H23J10ng75xEJeMKB+ZeIcKSa6+dxezgSGEdMIRmx3m0GaT60IadB
Ig/cye0CP1V4yH7BB4Z1yiRrgbyGopYZgkGWzJp+b07TFM7fAtgbL11yi1ofU1BmkkDqdPjarYTU
jNbFqbyBqDWH2bqz+0/mVEqfObIWn+v7S9I9CWU3xaodPRFs+BneqGZAychZShuB7cqBG/E1px4A
C0YQD3QJkBPLf4XCMFZGeXDxhprfauLXNfWfb74Z2gkcr7Y7d6dxFw+WEEyv/7l/d5xtgQMZZ41K
+wu0dgHFHuZVyWb9DGo08w+JE62Ry10/vwsJqo+BZtcE8EFOKgv5iUJy+9YcoHoFqHhjVFAs1xR3
7AE24BcjiWQ8hxSCDKDZF7G+2o0q5e+Cc0zOU6ocKooCCumiSyWKck671UXqu4v3U7DiLJlUbNWN
mKfyBTLf9WKLrorL6qIf9NfdiMUYL813W30owTU98Fnsfs5GZtmeaZd4/czvYrZ5y53N0Ab8Oulh
IxwNXQShMk8v75zEweKEPZCnsU5KSKyw6OTNvndNSRpvAJrrwotlHvNa2r2QTYg5G4LXN2XISVC1
2td2uRAL6dIlr974yI1FdW11J73GiEYgaNHGJlcSSWOcqJkO3cxp0Pu0Dn0HNgPmtB+Cz5RrSD1Q
HpRzEjfVqpK0At0Eri1C532nRQBGAiE3u759QZqT0lk1ueSBJIt4NGpZ4UED2w97mpHHN9w8p3m3
xgprhk6bOQSsks7n7LD0y9q8+5WHqTkCYBO+G/BPP2msq+M7cbaPCiO5eWXvsHY/Tj5AZryEo+5a
+dg5Hpx5f/2il7ZbUQUpZ7t628ysgnHzsQM0E8kD5WA7gD+2KchqjUxITDtp0dlimvX42gpLeu1s
c48UPt/NjBSwOwzQ+juItUTipji2LUsrCqnSAO12tMt29jxtgK7vkupvIVRcKfavnWgG6Or20gON
EEK6xV2ScHmWqatM+Fx6BXvyQhammBd/vtAypv/8S7g+TA9xboEXYseRhq1KKVTmUVwXIJQeUuPG
A+1W30trijkr2gr5I46pdRFcpWujNl+5srHTxFLIZCwJhQ8r4sGWI8RpBwffeRdyYVPNWJkdHu1m
VE68y0MBH/2w5BDwiRpQk7DSIcAkrtQsiI5e1wh4bR/XnoERvbjl3vqO7OmTgGwf2zDeWio+RY/c
tH5avgoOlnojOqj3IXDusbYt83QqacaJ7nXfBt8LTuMYKvcJ/up0D1SAt0ZFgPs7wuuSLEAx8vZu
33jNyQF3CInmBPO2xT/AkSrH21lnLaHsY3ZZqfVrG+oqGqRHS5a8MZV7VYMwjs3eTWe2zjxGbwHc
sJgA5mL48y5UdYM+Q9o/4nHlK710IYt/ykqbvQvkganAmhGwLFuuOiFOARm0k6c2LktTgQY6Qd6O
uBLZvE8d4ix3NlevRxWKkeQXqkI6ufoeeZeDeyBWSAnAU2jwUhn2MlnOqKFNfFqUvgd/VLMsb4kP
X6Hd106Z808V4mQJX6cXAGKfOYZtwih1K4+G4nNhpc9VuFVqApPQIksyil4YW8Z1vvX+7b2RQoBX
OzicumghKmrFQpq1VxBTugZ4koF592NEc4ORHniz0eaPJajEjYzXjdShnbZNL/5L1xeq2PXxhBvi
LynjiHaq9ql/+1xXiC+lLfV9syVykIJxtNvmTU1c5OlRVkSEHTzJe3zZmw80Ds+abceCh1pXDr4Q
Vlt49K2tQ3aZAaRmkharfxic+YOLEfZ6aNfeosMBOsM5azs4wpqTBxS0l6tbNf5SyBGbLoCI4vaO
2Uo8+xTEI7zxQgBdr/i0BTe+rNxSHjHriZhr/IOQ0dG32K9SO3CgnugbRJtg/R1cVcpC/5pyTQr8
ISpO24QGKnZBbGt0GU/6ESJIoXVrTYLOq/RrsW3kxQo7SLKCivY/jQkKLK+wv1wU9TGhfEP1D4tE
VT3zc2KDD6YWvGUHO8W8KmNXuill9a8H605M4cP+IB2eYce9VRR8XNrQxHqyxvmuzXy1rIZF9ltM
0mb5/rbUcCTWHO5Jv9BnkldB6VqTltuEy699oc4ZI795WtHeqOfcNzVJOPpmurlGZjzDKq5h8II1
UylCbKCbcSbecvgdwgHa4Z8IK/Yrfd0befwxB5h1zjmtjcgeGCYgex0sZh+wL+/7M81eNncxnw+y
UyJ5/i91qRXGdEbIZiAakMDZ7M1K7eWdPpkkBeIz+n7LVtgtlYypsFeRrUIFyTs0U+MHGh8PaQgd
d4ZxRBlBT+GgMPvIMwP7EzuqNvR7k7Rgjb3Ad29Rjvye3JJG+PE6hnRy7xcCd7uW9H5j4beGO81L
shpkLfEKP+wkwqbAux25aNOE3H6BO5+TOxuNKCiPn7amddULg/EaCAAAHk4Y7VAhPHptZ8VDRfxW
8FszvVSYmU3e/IfyUaq5BtyJaFgTqjlvUxsccb01/6ZHmt0qY1gk+ZSgwglZma2yqGozJnZIjh/c
zokAy6pC1CBDaMP39MSBOtUptGD240J76NohK9Czsg+edS/6GMlGKXGOo7a+dze8L/wxZ04o8CIU
r3JRZRYiEltH+3x+rvJ8EZUR/A0Js6PMnNxvxDgfiK2d3e57Zl3r9OGr8rkCo3DvTB+MrFxkZ88z
qaAv4rNbygk3P6fXA6uJJrbyBD8mmM3T5HIiPxovythQA22t5bE9Po4pRiXHb4LZqpHjloMTKkgW
uVVaUmgUqg6rGZ1LhdbvZibNh+Panja+xhYfSoArZ7zx2JiJHgbSzTlPN53nrlgayf3ocIJNA7Yg
iILWREo8psqrGeQjab+Pnl4bBciVOB06olG+XdcLrvcDZSBlLxKWWhlx8+ztZhMPRwLwkQGNGDw9
badWMzLvIYxRXdahEYvhZsf2o24XfNhDxNy13jT1d6kfFq6OEcIELGgwdBhAWN9xh8gAkY6+f8HP
BNWUvkHKT+I2R4j+YEwvSLcKJiC4szCY+WaXsjZrq+BMQ6I8JgGCXwC1AeNAw9m+QwdqzOoV3Dyc
7yTqQIGXm/w/32UivHqdqEB7TB3DPKDvtRB/lN2vdLNEr6w2D06xFF4VLlbPnbB7K+ytO45DjtL5
AunHUVBW4i5dLhJ+jDrcA0urwjnxxNx5zHZGIenJ9m5MnfmED8/ZOYzjCp+sAZsBDnoI2e/gMjFp
W4J4raE7wNtMr6JPGszFgGMepFQ/0ZK/T3dfrvWJ01HwHycckcYoauaC80Xz2Lc61czdow51Qwtv
/M+yf5rFBHfKrdG+MP4je0oOs6o/Veum8z7/+yqwvQc7IcWnl/bFiZ7Mk9K7OKBaP1Naot8iMTRw
pGlUDmH4Xf4zT47M/PtnEl5GY3KNiI0jM6quSEW+jY9ERRlCn4qmrfV/8K+H22mew7u9hdSiszwl
wfXF3SGHrWZCov6cKUeIPOsnYJBtgkaMc7gSY/ICNjYi91R8yMsWxQ/2F3NxfNBzMFQd6meS9reA
fUcdgE8LUbqZjurYTNjGu8Rmb/qpeIOazLsKvwz7CUtNGWEwc2J7+JKBxSdhvYwc/CuzIeXhki5v
gsgOYGkPR9Hc5uSx+5YeXkkxl8ztVy0//I2ptXhu2f1X57SDii6y1qXhYDJ+A9eaMMQ7c52a9XfO
7/fg1+Vg8vSduckyJybQcLezhQnwPmGDmg19cPREsRYOQ0mrJsrR+A7PsfRh4oKVpF6RDwMbuRQ6
JCXL+2LpNg3pTAWyqh9umMHmvl3KsoBo4oiBXDYPzHAZ8JJbuRRehLhf6Zz0S1kCW7KbVi4l2nrq
z0sgVhrAIC+TwMBXFNHq5lJetCumXxxoTQi7MdckM5HyXoiIUxKaTeAsPgG7AXD7+1nDAlFhxgRc
pq2PmVMZ34U2nefqUniIj0l9FCOQsXIbGOILXcZ6xFy1vtLvATCdcdsAhUxLEg7gTuOG3tQOEuUj
cRwWNnqI/8LEglXD3BJeMCc3HEUIcUcSxmjgtNejkDNU2CWbBpfMaOVZAM6fDrUN18wZPKYXjN3k
P+Gn8f0OA0SCxvfGbrkTuO3jSLoa6on9Udb0UWLCs86hjOdJ5vgFjNeSnKLDR+vF+u5PA5RHFMqL
CAddzt853NtKt0Euu1k/hev7SVqV3fLRTX5uT5vWeNqacB20HQ/vjVIcR0XTazdKbu6BUoKTtvqW
SuKYFLUYAMh+lUSD6he9M/aSRd7w/9J+yTQS4wV24vmG17WCB5QXz8I0nGz4HNQJUugc5m/WeCYd
5xhWOTx8e+RkrKbLlRidxJ4fYuwmdVKkFyikh60glrspS5bE5jquCbx8K3sSoLUwzmSm6zXyqDqU
S5KEN2m2TGUQemHkJts8bYR2BJ62269NFBr47G3Xm9W7hgsnve7Zmb6cP8ZLW4USKZgEH5xJgEB/
N/QbbzgvcOD7Rtfd/6ueEMyFi4b7OUEghg32flCOF6qbESW4XYO1mQN/0+ykWRbYqiwha4S14vst
LjDi125SRNLSDKC+Gjl4g71sYz0/hHnW8SOvn6gEvprv4HAyqKbfnzaSsXociUS5ZIBKetb1ALg0
uXor0vE3qVL/FNX42Ehj1fXt02tOzy4ncRjG+btUsvbFIDJ2lH5aYtcwq6GNdZp2xNdiC3ND2ZNx
eEdqyOqRswHWcryNgsvDii1SBr00q1jTxEn6TEmq0exwyfWaKmIazz7qJ7I2Yc+rPvNLKe9HmKmb
PvKGQ7lrCjIsm0L9oqiMHf9FQaDH2IjQdxxIux5EasLW2nP2C2ywbCljIDuXCdLreUd6p2Xah38W
/tEJ5guArjNwsFRFdmCA/D0nDbUfVI1NRBnne2uZnMxh2wQznmaK4FGFAccZ7zuul+llFntRiBwf
cnim6OKcD+Gj1rksVWm3zAjEu2yAG7l0gy/f1JqNiQ/Nv4mXVxCemw9F6vjjbtAUpusf8nGQKf6D
GCppKfzQCBvOqS4ZR93fz0DeI0YmXv3Sh8lnGbl0+xn7HvXU8/Nh81G3Ts/GFS/6DTzCGums6bQq
MlEiauiGE5/BQnfQqlSkY4hDYvxb4Sov2j/3O3s66wjZSoT/z0fUvr2M3kKsRgjjeIuLLe2ADk08
SxiYKN+idVh7qZfTQUda/EaEEuyfVwQiF559UExMXmq27uMskWF50hW90dj2JSusNNxGffLqOG+a
8U1NJwEA2/Ois80xBklyMjEfVCcBJUO1Xc/idVCItNgt/wy2Xe2L+42N3d8VJEdljpzfyo1zbQTm
8odGgx7T/U25yeP2GIBcBQSAIG5VeXlkPYrwyTIdGYRhvgO9OF6U574dWsZuBB/14fpDIKG8bVzA
xFcVt7WXe1zH7bhaGHA3mk6zo62NHB81hXeAbLaJzJzwuQIdsHL620xnbKo6pIdRwzhRo3Cd5y0B
ZydlzauO2YyTOcINfoKL0XcwzTJwmRX24zIZs2nE8k/xqBlXOVjgcUlo5SknR03tHJuZhBABjcMz
uc6XSRnDTI0MXHUW/H+NR4CrVWamVbiUX7v0nsamTAmHvOhoy/W+0YHTDiJtUe+JowO/PqDUTz5x
WTTqU9u0iX2b8fVwxkbvMr+hQGgVsxni3+wv+Zv0MeRYyvw3+dlWW1ryLwIr6qhWA3nNCIqzMJCJ
b+wRWBPXAUjoNzCXfHoGtzsqoiJ1P7/OWXFeI17EB9viSydLrOx3Ms7BFQQ7oRGuiKvzw+CzfUNq
sP3aWM6sJbknAo9CRkU64cywQkgRfRfVtnEz667iQSYU7Qjp7feUS8AUZxadJBsE0RDk6cI6fYY9
RIMkVhWxNxfyYihI77HWRVGUSGgouetfymJ0/AevgFbGgAu3n33Tua4yxUhgqtXFZKifTDixnPrD
F/lrrMvLE3Axaow4/SE6NeOylp0zagFi8vAPB3hQcW6AhwwwbMbeJyA5PkjnTPU8YBVcENzp9Tyz
WyqF9n3xe3ygX5+In0c/RW3p6zU1sCWpQoF4DU5ghxF1J53jGnWqHX0aWzkWvm4fF4azqUwKOhdJ
2i8H30e7ZUb+/QMTSIv5qLtJeLu/8BN3ivyZXuvBuR/dTf0SToSwVp6rSC2aSMXs99ay6ho/eJR5
4fkdjBYY14kc3co/dejlkbWpDzQ0IebETmq+uROgOsEX6HlhZioPvKbtKx4JaRWqm3SRh4YBBKCS
lqie5t4q6xvxI5znFM0sn8MZgX+S641wyAhK5ppOHRdGwZ9J3XvmquGxUcFrDj+ZLnqP5F0KH7+K
+t2sMse54pH/EqQrFxJaNpl40u90afLmSWlg7xIIJEIFNodV1JvBYyPPb77bM2RorQSHF1CN3xPn
tjrDKXciJZmmIorDcvu+S06wtwhBWSYJA4smLK1RitHxI8Csvqk1SHvLthbTmLgGvOYqBVayX67H
BcTEE2ETnGWutre2n7ma+HyOaubrAXTWXB8KixqC6S42WLto0GpIrEJLpSmF26Bduo3ic5p9MJu1
nEKlbCiuWjoITLfI/YuxNKL1+TFNJoP5d6MMyJfZ/AY2L9OKu/cK2aB5hIKg+HBRQ676YdY+12e6
tP9fHaKCRA0gxgVQas4KyF3Ff1CwiQxbiusA1JzdWsMKg55vHMIjS/ZGCAeGXtBiX038w4Rs9L48
/9X9f06E63JfnyMS252Z2A+Ittjte58VyTAV5nt147wWCDHIIn2x8JoOb64K7pcyWaIciMkkMCh/
I4wg9UjN0Zhg/LG6VNAl2TtlrYM/nOR1Lo+9cKvtWYNJSKYipGRzDR9YpJTiO4rncaG+dNbnzs59
tBDqJeoIMhkL0hgNsjjmFSgIiPLj6Y3yf+8h+lxSwiN+XEVieKbqsI2qjDgu+0kKeLOCD9IdhEnl
MacN0PQ6UDFjGyYPQb9Ouv5eaU/QJYPsLQfm3FVIedrlZJY9k9OJISa7EaQ6zjac4OBrP6IcOgJz
sfPAMy8/H+4gFPO7MoI0v+CB9ropSYbuhTi17mYTKMsp8VpibZ0rW6MUhqgWOkEr+SAZQ7cwQlxA
tNM7i4jYqaZY6g/HBGNpBBetmqKpP8GEcQrtd24cVnZQLK85WpPLCRZSFbkX4/SU0/kQc54jqqYZ
qFQtDpb3tvzVSddnyK9Oxc6qFAIJ4EB4KiBoKz3grz82JjKfTjrcueC2ge0sGbvbhiyz06O8rnkN
XaecI+0Mfgywq7YhmhWzTuv+P/OolUwfi9qtVzp1M14SKxx1LEvrdB5c4wk9OSj2VhzxL/hp8h1C
XXB3MTzFEfFxuvt7K1cvC0zBMDlqoFXnciUQb6B7GXMjj/B/0hRUOaxx1SkrPws5h7Poktqw9Id7
KqzjX9GkcRr5phUjFPxpmLbeKFjSQdJFPY6G+I/j1GN//Fv/xFFd2CAe0q17XUdNfy6b4+XIgh2D
UmQLC6ivSBCIfVyTCLT/Z1I4XVCiU//N+ujR7Jb4KvuymhtU5z+iRX2PB5fSQKhAnYrM7c0Ko5rR
JeXVn0612KfPwXVHdcHzBGdgYSxTJBTJPChbolhiqKDpVcsE4BjqjwtxR0L6Hn/f3fhwJyxk1qbI
uxaKeCT4LIHc79e3vA+4nCMneMasN4WBH9pCb8c4YR/XQ0qllxDPHh1KWlc4QLem4sJ7dpmxqXzt
iAmOqIYSI/J7/RfDQt7B30Ug/XQldOqYc58moZlpe/rh1J8F6F7h9qCvNi/vpA4t5Q7sYEJlJwsN
AbAXwCtohfJWlqu804P9OXOPRrv8HgdpQ3EL6aWWD2X0Fw31liE3v1e5hgui0oyc13WbjE7MEeFd
oYc3sG7FwwFyEJQDtyZIuzV483dNHEaCpOOOkVQateCVzvCuTer3c53RB+Je5HSs7vGC3iPWejp/
75/4M7WaEut0AFYQdZyTrnoCXytar9HZdrMtmJbmLc9pweu3YJ5UA7Wfkm11dJ48nhDEhSsIufQw
+URl6BqFgimnQpruzoRRXdAf1XQa9l4gdv3yEFmBaQhzzoLJnDpmV5TgtszSArE0PKuPdJ4gz6Ox
6Z4jTIzfPYvlvblY7CAukZBtBctO0J6ckyOA0MYDocm1HT9adiDCWXFQVTyM0Cz0xLhcyWCZulYi
rTz5l1ZjtucuD1vYkajCDOle2ooVNGQIyCV648/6vpzuuN8Yi4/1Ha6m9QM+GnrBVXoYridtIzP5
6rPH1VBd+X9GXZprsfbgm97CAHagttXq+lqloi6JHy65HuG7NH0sGV5tjGDgGmIekkXLDSdvrxDx
EIA6WGgtScwbenrBDUFf86nfif46tDMRiwhVa4+ZdyXCWskobYiupau+ET009NUc6no4Kc8RaoQt
HWiWeb/yR1QSXuFCWGe6EjaDsbRXMvqeZUSON+VZhuilrRFdFuRg1QlL0W/TqVKlfhbExHDNw5Up
UdHimxY6vU5fkNxsOf1QdLTPnLTE+OwX4jIns+OlVpX2CLVbq1yjawXcgdQcSOREjX3viqkgkX4O
a9q7as3LezRyRlx8q5mX9ocR1ZCxRPm7H1rA4n0uqkQfTlUPTO2MT2nLJnKU+qq/
`pragma protect end_protected
