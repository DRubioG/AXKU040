`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
HfsJrmGIL163EJ1QN2P8dPrkZHUc1GN3XrOt2B1bnGZ22+1gIBPPzCsebrH1Vj2c7zQ0iP7qjSOl
hQEpDzVilQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VwxwSsaGBSmtEHiQ0wqacBF0mrqKArSeZYwc+YJyKb+a+QCkBmztKcYNXRK+oQyKfLdQh3JPy2SR
JxL/qY50hV2D2W9zsvrnXpBLICtFhw+DwcqoON5Gi+WIjMXPrwDsiJZ3hV9ztt3eAXS7Rc1BDf/Y
41xGu3gJXOf4Dr70cRo=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KYVEd3us7rwB7ABq5Jrq922AZ0Ujt7rmmXL7/niiTOhVRz0f3ENmGm/3ZDuUI/1F20STyO0qKIKB
mBWyNC4li2ovQwoS0hrUqLsz9YLUtyU9Ph1vUsCFsnfb24FXjTzbKIREGk0Rl6kzsahR43A0LHpa
pWkWaQUbTPz6eImAN6E06pYsFHpKweASTSpfR/pVdcAR7QTNvfHZPtqK1LUIL44CMlH2uLhhzchT
5bs2g2U9x1RUQAyllVeNuHuTxfAvO/jRlAhC5KBldBlhlAZF4mLI2dglyIbBaZO9UYwvd9Jj0olk
PLNlZAWJaeVMKqEwJ7tw8xPTPI8qsQNyw4UHbA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H/dAtRciYNV8xKTfomfS0t/4JNfnVr/ZvAuUc51kX0e4e/WY3omnqMt6T/OGtfYerKDqenKfGylR
N2hjYTQCuDc1O2DyoEBJAgRJAdkoHDqINfngzxnCOayHooiwAsUTxVGoIfcEYr51Y8ogZHHp88Ae
otXE+4pOMe4fW4IBf1k2Ztrjoy91sTVzRVZAYFZHDDkcj9PBRCFlV1jGzaXjm7HobZwlNHU1tIEv
y+S6gh08UhSxlC1e7LQUJR9crn4KLl2AbyI8HBQC9ZgWWyUolgYiOnRj0NmEarPqOg7FX7yYrv3L
Tvp9b5BYHEgYi65aeOUNOMcuX0vo6hGFjUU2FA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FZH/F9v4Cm8qEiwNJbjqMu1aB99CdzNh562182N7AJU6ZeCK6T4kxzSGD639e/6f6g7JoDxIbyid
KzFPHuI0eRG/Sp7XlJSuB9RtBBBxJ7016JmP7n9ewttAsIggpmOEvRqJrl5PVxQ38H+2nOxyzAmE
idSiOJXEl2Lg/ZeJBbc05OV5mqhmNg3t44chTbRvz60+qt19bylSeJoQ6huO+nZHMkgxWsiaMM4T
P/bEfW4unJwvYE3a2XqwWmqOVTTSahBz47owqL728cOKlcjWFpnNFSmoctmAdFZ36ZbeT53mSV7y
lbzF8ANRHiLj37VdI6hHnibK2Tzkcv9BUGxh+g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GgpabFefzr9N27bmXpx81TybAeFHtFatepnf52KMEAkx2SNXtHvDQ7YRODzUCba6nOM6rppHWR22
hkpPiLPCcsHqnjhWr2T5QrHDZPcuWybDBsh8Ox3HspwWHYfAERCqeJoFr+juoqSlqTBVXi6QN9P4
hwrljlSNApHD+eMtBJ8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gxH7eGu4ckovMReDNzzRxQRAwfGP633VLtDpIuCrZwKocNGopmlPkCPB5pnebWZdal5JZ6CoWJem
iTuwlYOMXQkpEE48b5P8cbEXjj6ImAKWj8TmEZOebr1Xo7G3mALxQzZ0yweVhixbfz1pk1E6WvbF
o+YvWhNb9eTyv1WEdaY092cQjpzKQLg4V/rkvUZ0SZ0EXZh1pFnkUf9jrGK5mriNLN39eCCT5eJp
HWQu952RXCbONJ6uGxtHV/80LfIuonuneCAtSkyN0u+ToxJMWL16AsgqQGrcMDtNCJN6igfEFw4c
hU/FON+SfZqfeQz9IPz2igQ9efgZHZ9dgtVPwA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
AVQCIWAosAAfom+rEErKQv3v+IuwG2INN/iyfccwbAfWgRCcwBOd1O+phehJxnbFoBdEzf3XaA8y
0ObhXficiu0TarMQvoCmxb0HUP2fas/zuBBXKuF8h3PpWhbyJ7Eu+iMX0BGE3U7Kzn1eIzGD6Sns
GShYoXTzWrClpW+vjuyRFdz6Z9qGj5x+WZJ0Wy8Pbs4H4L+tYn4Mt8nDrFQctnjw+qPPt3rZHPUU
v+RqhsoeAVl8OmleQMD+lljZcHMzlHteUOPghhgCkE4gYrl8c7DKFtGPq6lfltO8mZkmHCS1ko+j
pRvriNDL390PnswoczzL3Y0GsasZFA2nbaaxkjqBegykPnroNHb7KNAPECgKVNN0ZSppD8r3DAs6
vcJ170AOiKcPiwVnXoEnFbURFAuIzezdvWKz/Lu6w9IHdk5nx08B6Kp8XY5BV6Z6GYfcqX8Ja8li
7PYZblg5SyqWGzGRnbBtiBKIDPSqVf/Q7E/EvqHQKz7/q++nYgZisjZ4OweDMu0uG9mRzdehFs4h
Tj8dA+d7lD10PnOS7gDHoF8FxNBfjIAk0TR0Zac7bL2R9cR76P7SpCvp+NHTy5Bg/0kaLW1xzprf
VDgQpiQHqDssxdpGBKFlUtYIlLQerjirB2jZA2ZNNEys4zD/mjAbYrd+PBvQgDWvEuybBA8RkHEd
unAc6sz1Yf1U1qKyqiGXYX6RUjc8cHne1nlbMREmFgJngGtgpx1uFXdQYbhgkro0KbQtQZdf7jEH
KXWjgyCkcIuU6lSsr3tVRfHCn9ATsUpvT7ovApXdIqHofhEjfc/Ko27SdTa9ChqTP35swhuZgH+8
hNEwRJieuWJZEohvxfppOdY48lCTi2uIN+DnHq6IYV9YtPQnlFRb/LvlXQQ3c8Z0qxDISclojxmk
UyV9gvnkLqpX09bIjloLBeGskzfhFwde8mswIdCYbNU/2MvMxWeMCOX01ma8QeqKCYi2D6+dFRsf
xeO0z1D4dwFlTzism68+xnNzJeEeSxQrXq7+zDPjngTlDjpD5jQkeOI3kb3ceudzgIgtj4wTdHjN
QSRfx5lBKvDO+zBl4YXZ6s7IsnpY0n/EEfOAGnIo90d875y6P2Evg/XTjffjgbDzXY99YZg8ZDcH
+hg6aRV9soMxAyJA/+tYouxw0IkZJQrC0ttDVV0+Zi+HpA4lNB1Ope/QxeMTbs2n9uCHUVuifqMN
j3iS2xEP0qCrioYzc8jepZmjISNYN0PPf5zLhGG4szlHTITv8+nxNxJJs6ruNG6JriTdpepwBlSB
yRM+IksqakGQQizdKxBf+a4nGWUaA4zkSGD5gIQIGWqTbeB/tF5C0XqKbPKi4zGfgsX3btvAS5o5
tdNB5rWVZwaenCsSzyFTGupHDweWFWpix4g54R1WQDU9SWLFxnsiMRcqQqoWa1M7MI6wV3kciR8D
TwGBDoTDWf2ogSCarJ6P1xwBEBgJFtk9smEA98tTuXeGtcX3JKGwpk8ExPUuPMq5xtTKQ25PcZ2J
0/6uhrSTD606XQMJyIuEHwKGN5z/vgQPHjhYWVNaes7RTVmmdtdQhAQfByrJirbd1VKIp0ApMxQf
fsfw+s8zFuSTSK6KkcpALLQU9lGfCPBLn9ynDhiYX5FEs62UubmL5Qq0KISen4DadzGzZRxOzuGp
RBeA1usrSnKMO99cB3X36jzkgZxc1I5XaJbwAZmP1D9RzqpoFjPc86FX4meJWUvvkYedZySpbgjs
vaA+UKMTnkRYHIvjvdzf5jX4n8XH22sJnONFTI34Kj/DfU6FHzhzIl3DQD1xHIwx6KfCsDwGu3tv
UAgO6KqQ52Xoiy/TrQ8/eKgVdEWp3yTdTid1uFBCWBjdeFMTNMUeJ/FZWWIjuAoJpbSDJE5F4UbE
PfEmQTWTgBMQT4kMIzEyexkyE0wLnP3YTbpZA5d1q0U7iGXJU6CVxdLYloZwJXUTzo4UOV/lpz/n
1SX96pFLqk+yayttLexYdfOp3+t+2z1AYByQ6iVgJncdooEQUv0Knoyh3LcSQ/NqFUnmKo3btv9O
Ai2GhFobDgiT24iLvwNdkRUcAVcJ0DjbRmAuqfpnt4NtRFVkPpUn/PKgftTXOizW5UoO2UR+D95i
Gzmb3bCdogSUNYc2hXvUnzanJ1TW4Mvcv+cYH3EYS8p7T4OqNwAra+t/ZYRc1RuwvTcy5y/LZhuu
AVeBqL9GRwxqv3xbf35WnGogGTims9wI7O/RVTjNTfdCwchr2zN/WU3EVq2qXyaIswb4w+PJU8tD
3mtSOqoybqQhLiIw9Pok7of/ImSvy6V31ty80f/roKKG8Vj96kKtniroSp7piXQKDWwstP46I8S4
KccxUn86kjcSpYRLAnV8VfNmtgTXV5R+pBlF8sJBQXiWBojwZcXv8kL/7IDi2zkIMNeot6r0B9Uq
Aw759ahrZyyTmk5fUzzI6MDe3vHwhCMnpMdhJ3WrAq3kRQJaPkDTYXIqThkhDPWhoan6mjFFeZV0
KC21JQZBT9BIV5moagziV0Ou5cGfR7uAllA4rmfWZNCpWh7fdd67bLTVLFKyUfIwxXvhiyvDNLVX
i6I8VdXFAwy/SQ5vClEVTlbJgvBih79MFt7VdZGUjFFWNirGhOTzY0OerAwwDZVs3QRhUd5QWp+V
gGoms4gHngKvvwr07NnOcjyPqupJkZ3+ZIubXo4BopzLjq662YRb6iuAyOH5RLVKwCvpMuTym7z9
Se+NAe1qasuWnpSqUROyhRzSy0mEDVdgvMbkr7DtUNPkohD+ylikbSDB5bttOaORdrl8bGSaMgXh
h1um3XM+T2VatD9cfSZSRPwLTIu/sqpIU2Tl7Qf1wfttcwCWCf0Tnf5FI0VXSgAqIk1DHLCRejWR
U+SmiHkAcKiwzNsVtMy3ajDEkrmADUb42dAh1SboKI+tBSz/yfQ+Qp3MQDy88V2UyFEWpygj8Mol
szczJL7MMgtqK/RggRxPAe84jiRgaDjR5csOJeyh7batR9xCLKKbBcASCq+mlilbo7pqjwKlpFwC
NlfzJE0pfmvdciQweJMeS5Fv63DXkDzIFiVWpMzbMsHAz/dpwyux7DmEPjH+U/DgbFQqraXtjmTO
2QYpg6SSDCXUmxS0oKhLIpLbEIGOuVFTAH9vkhkC+feaPzP5/xd2B5CS15jwjZtxGyyqQsudwOuZ
/WiBlDaxVw6MVHYzgCNbLlDNLJ1eAqnuRDZHhJu4YZQ44wiKb08McxwI0JCxUxtprpdjJlYYv7RR
e9gRlBHoBWy1Ak+cq9s5HIVmY4G96ELXCFADnkB7ls2IBX1P1lymmYUgDmOQXXXWe5Bg79BPMV4V
UYIg5fr/MSlQl+J8LEzuibs7Otg5x+Q4Z755QbIMAhpM2UGfsldqVJypzaxp0j/fiPTTOFkm7HK6
ObD/F2BrE4je4bIJyY8MH5hOlUSUWj6c1O0s3NVB1P0B+tPSAfFt3OUrLwp65EiMbNGJJWX+JEtA
4hU1SEQusSZTKsNyjjFqHf5rYFofUXns68np2pJkBFTDoTZo7WEqWKwy0KY1ILgKO8qdlFER6/mA
QJn7buILkNMMqRIib3usxwXDlwCfc8Aci+fKDLDVdnW8QD7KAV5/yzBexREzlZFS0ZrPp4xRc5jU
mqy2CKf7mwrBPKxId6F5q9eQPzHqBkYV7TTLwMUOI1bRoJFWwr5QQfLELXXUoloq8/Bd7xLUS7Hr
YPC84YyKEePwQvJrv/bXKiP2+ryX4irEwxW2ZDINba+kOFbKSkaT46cxc7MMb7YMa0KYx1UDK7uk
OTDgdWURpW1YRu213H0XyIdZB05PO941arDtNWHhwDmIeEC/JaMBWzg9yr36P1umUMWU51INJ532
dGczm3thYZ9L4oHaF9gbmBrWVezAkqsHW6oiK+gNn6+LGMnqyzIjZJ7RePgkqMQ9Ix7KgTqLMP8a
I61IgYapaVA8NiDpIptG0CdjbCcZLkd5iRvzc19nD4IT1r8Q9riquuZpmDc2Tpe16uYBZ9Kb7dOb
FiDK9dd6WsT97RZElfa1K9fw/d808bGxy4j6EXq+WbdmuakYX97UzzIJ7FOZZEWtf/A7a2cJmWZz
hCYi4le47kmooqrD53t/Gt/YiKhtGkymZU09ocWp9GI90YAA3w3Oex9PDJG+uyTqjseFF6aD34Qa
lpQe4/Nd+DAr/QFLTMoLkZ9KmFrB1j512LU1qiKMYDeZtw+SEV3AzkTF2JO+6q59tGGA6uxLIkoc
9betyT2c9pYR2yYTEn+sgIYhgPXLK2ysRRA4xE4lta5azT1NemH+YqsvJN5ROCudX4HcquHOlPS5
ROuZP++M5DNhvG0yH4m5TGtJUZ/F0WiopH1WQVWo9+DdhR9bkSZTgbj8RWSfV8tsBrMovaU+J7Ce
sE9IQokzAUx7m9YrQNImeOtEGMVzdOktvRPx7lLk/8zJTS11PVF2NHbqfTJYuQDwvGp9jPWiye3L
2sQmrgVYbtiXOwivNo/pmxO5TTntL+8AFzoF9wuSJL8I8OGtom6PYnIjJcb37M5JBYPkarIvrc/i
TPmhuxZiuUPv9cT6X0hme3XGyvWNXsXQPct3mF9RFECxug5QGDX3Cb/SqnlxHKcRHsocVq7CCzQa
Bdy5CcmH0paxcpNhqWhBfjpgQo3qMjFU0tAbTnk6Q9dtuRHZksjo/vSc/blKvHQ3zgvyv2mjb31D
5mP8aKToeZAmpe3Ny8VvGIbHjUTe7baa0DKoeHkpXS3q20E8sdwMZOQVMYP08gu5esm9lFXYKrlr
glDPs9CbmDa/IEu+HWBS2nryvPs2Prddn2K6c6k/Z2KPvPNYVH/F9nmQomjuYFc5O51wVEN1oBoD
wQwHnzOmtR8WtnfPl5f3iDZnhQUCKrarXDJDqBV+MlnaEFMHFKVHFIoyvDT4H88ORIryqampAH4s
GYYaL3QF1aL9+gjnrsL2mIHvd8GkNU3+m0gi1JwWM4Bw+PJb1ndpaILmpLXZ/Kg7k/YRcKv04349
LOL5D1K9ZpBhlctCxM4S/lkKN1SDyhS9TM2VQZQOgCE3AUUFn/cRlyoGgtPRPOETE/BldOlke5N/
U+9w72TAvxHDHiFEFp5Pk20+LSWMVPC9eYwqgjmm9Wm2GAyVJvyQhI2oxY8TNHeZXljniLTKNLS3
IkgB+NEt7ArCxVYN/DhYTu1mh8JMok027No0aZVdXb1LlCrLnS03S2OC6ZgRVV5DRQlYusZz8gQY
Lkl9w5MrC76LkcsgqU6YWBP0E0PAwypLAaie4yrblbxNioj5LngnbJbzb76RNSQh2yQshk1G+XjK
kkosDX5w4bGWQ82icCNL9xQVMPnm5o/utdwltUKZGYLwlJDlvT0k9vcBQVhOxMtZhrjEWVpHU6CI
ZwOte2XAOQTm33pbUKPehDDmQOB5CBYkKunY5RNDa0dt4pATNDkm+JyXXEIAvjNvAdoR3qy7tBvz
612vDyDf84HGZne5yxNbUWbsTzD6/6ZGyKrKB0sf6v8wdn7OSAhjLholtLGzsHz5kKfENzvTByag
f8gMRuW8PHP+YjFMZH9bY3CZ1W0vfxVrRcEBo/MwtvhoODvDrIWJ8xAjwFo7eFS44+4Xc6vO8Dsl
JEomJsMlh2cguq58CQVoLxmMVLLhPiPg2fhbC1+xThLgMYfxM3ytG+EG3wdmymumR3OvuC3e1Yo/
3vc7p3ChyvCNZinv6TJGagnK8ZqilDVBTz2UOJrb3/buLtXJC+s0s31FdfwNuOvwode3ONaFTN4f
13/veE7O6AUfBvoSEbQC6WE4LfgjvLViCtcRYNrwwzitI3RChoKO55skx9nxGbt6gxRXXX6dlMI4
6CyKaQ9MHTeHMWZBHd77O4Wf7me61m5O3jcsLK4P89uBIjPbSG7ZSaddDfpmtlqp9lfb8M6Geokb
oHcCGECTGyCPgZrmLZLAipiMg4Qpk1bPTEUQHC7IrNusAIiNvWHvw3Jq/I1JlPifHOtAdPXM36en
S1Y7lCDnzanDqxWweWiR74QUPpRC1Q7R/l0HnEVIGxzNuSblqW2y0PEA6DnDGgZ9ZU+wfWwr4dOO
L19/q53a/ecS/5mc/bS4dsmGAp8UgH4/ndVpO0dCq5Ld6rAin1GzSEUhDrnhH8bVOncxMTAItvvd
g5HKhuF3ZUgSSDcPh9Arj2HBE11u7Oz326FnU3SK5YFDpP+f8iOc9yrLns2I2CcU2pb2BjMTrDCO
hpysAwYvquh8Ti1erEjszGYKLIvuJtZJ/PyD+u5P7MDJJiTVs635+mmeoXX38pQanLtpPrqmDOUN
oI3tOVTUb/19GoFiFeKA+kRSXhKfp79rRc8WzXRa6h2pXO/qKgReVV8pEbOz3ufZboyNnkot2y+H
MIFS5iffPfDNUDIXViYJrg+BmypvtgKldu2jushIEWDMvpDHrflXqoI/ovUx7XRNGkgDILKFJ/c3
Y2vz5MdLXwLpaHqbLrFen8sPGMwgykHLeVLk7+aKXpQSyyg6LjDWhX/ZC4xQ3H7Pul+TM76aWRlN
YofA0Q7DJbt/j+DopMALTVyS7Yx5ehJTuUqYZwyNE3Tl5MZ+zR/85GspRcXbGLRLh2OL07/nYo31
WJGgcQm84f4lTlmXsvy+DMehESL9gMWnAOEXKzfNs7g9gzXA9TMGP+52plwAAtqqS4Mrj4hUV7Ul
z7Q1VRU7vejq98EUVwm3cEcIDfsLHoze19fq1XELYmz5LNJ3khDmnrdY/M2Why+JbWAV+fvCG4Mz
lrekqsOsNbTjBC3kx5SgUcNWyXqh1DUUZMnkaMMvlo6cknnPXntstqyq6/iLPWCK9r6C1OxOvoRM
AufxMB5dPMhOw68xHk47BBLPiWV9+EgMxWV3Gvtl5bl+eaRAn3IDEprMeC7ls3/uKyFX/Ge6n8bT
uWYZ6b6W56dJtuW5Ls+UrjIxcYLad20deUNwri+fULmeqiQj8gMkKV8e1fxot8Sm+6/IcGH+NZ9r
0yZ865hQJE8NRiKEwDAaCsdTNUawqODMa+Yqqi1HFJeFT6GVz4jo7b+B2x6eJbLEbUGhS+cFwJC7
8wvHtGjjiQnGJUdBxmhd5bGtiooZORN39cT+Sv39yOqG3BOYcjxP2C3SDe/vdez38Uu/4NgQo5Pc
HAb4JUklzu1x9vWloTVdJg5a7AmzI9pVRrMUZsIxuSS2at1yMVaudb/Z1LHOqZEMzmq5xtBVU/De
vTXgsbDzNC9b/MjDCvRQoJldXgnZOJh5qIP/7gxglXGoi1lXxqZ9TvLeSmvih/T8vSluwcOv46hX
+AzVR3yOkVKl9Bl3CBrKhLXnrmUyU6BXv2mge46TgnJalovWZ8rByET+oIc/flhDXleCU7W1oZp7
i92Oz8vrOKDCZkRz7AqY7wLyND26/+Rsaz9OKRSYAwtVbXOzm8s2zjNPWcKnysFHcNudWXBhgi6t
qbxiMD0bvXKuKBXjLpe1gfj8tMn3tqhBBInKlf3g6p7SYEz5dJNw24vfD7HvxMpjwWpP7aD0VoYN
ysr9QQGRR/X+imNTY0OGnCwmPENq3Mow48TKLhVJ9uhGv7VjR5gnDqpfMAtEmTQxcZz5V6WgSdex
Kn4o/iy/MJpnPqQ1u9Qiq9OK5CZPCnRYyG0K1b8KcV3a/y408rdGdbFlLo4Gi8uZIBFFdamLjQOD
fW3MaBL6oxoBL4SbDI09Vuhn191kQMR4qi6wYHPMWjU++ZyZS9lj+wzyVKMz8+IrmwWvZkoZig9u
+EFht6bP51wdgffVrFU2v82KV7nOuccc1wBfMTORTjIUNVmxRQYiwNSM9qlc6LuUgxEOBUuW6Epk
pgfaBgVx3TFP2KTGlSPZgEtZo69vIzIsdMQ9zfx+kmfYXlODxjkWWQNnNABvnqW+wySJOMnbsa+Z
54VhV5+Pc22V9J2XthlGBCftuORKTV1ZyUTF6uz7ZWytSeTBKypEFdIWfzxzjW33N58B4GloBz2U
Wy83droCWKGXVv8RyfQRUwXw673lY78Ubje3zi6+8RgHbIrnaHlnw6FILCD/Ldq9wZBvPoYSbk3v
PqVL/LwS3uH9ltELR0M4vErGu/OuC4upSMSqbVp69yQdqQSDImI+jAaUnupwCAuUAFES/VDpyGoS
d/TDu5tgX4arFJvYic8ruYPrNuajfISGasxEWar6phAVWVelTfkIWx5IuClf6xz4jM+4WHkadHCF
Ph2Qh6EidDq3fTDYFpdy6c809vMghrFR7+I5tcZM3NHMyEIKAyZwa1Hwv0j5VF/KPO0pdcHtr/1U
djd20qasKHKNm6EsnDsIenayfI/hVpBLnVqvILHM1n3s1qy1SFBbkP/vXx/8ZHD9Fr8pYpHDc0j/
3xMN3G8PjQRrT8L03/CxTH5wixfOabVnUA9cMdxZhaYlPEMUO2s9785ifwH2tKKhxwzN28nRdcSu
LxeeazwQJ5e7ihr9vLU2wvaLDOJmGzj71o5SZLRInjRE628X5V6Y7CF2JZ8KXX4S5ORNeTjcRdyz
BCgDPKhNKfHdMUFlf8UpdLya+S0AxdViQaq/IhFrCKMEXU03VffFoOOk0a7i9Rv3mOKSsyJKb/G7
GmlF7G1uNEmn27HN4j+5s7dm9B2g9Jvn+cCVxFrFBTmuCQbHGcfFtjHPsXW8jJKuVrAe1jqIj489
la6GtUc06xpW4eqUxhVJwCe6J5afZgeUCvZcaa+gt5CeydCaEIG7BrcIwZLV/pN0fMURmF+n9TwS
qdhh2gY/9HWPPCO4RHWIUlKc7n6O2vJqHaHVBIc9aBn3UFRmZERqE2Zwudtz3I6TQR5WKbZ4/8v0
c7pmCVgNHjPZlj+QBHPbB1sl5kNLf7OhjmnInsZOO0nFQw2/P1YiKHgQwlhKVFOahmCv1LEJEgz6
LPgtiTmrGSN4sY7n4Sbdshl3UG7i5WRHmHJN44rEipKGXt8IVpJTVqx1fB++be00prQa2lyqyTwM
UxsxrRMM4+nxy+M//1c0uf1ROVK2HAoPOqWe0tOCH4mNry3JSvKCXzcMezm8Ef/mI+eAQCq3W5X0
e9bWKkhs/m8gYpbE0uGOwtkZ9vykC9jyYqXvfwxk+qCc8wrxW0r+xv57VnZ4E0+NPfkgtx7izoHM
m81wGqRve+3M8IBmB6QVQ+uLVAaYQOPOXmV4QZChzawXmjOp1QwI0mT5chIDqJpT4XWG75WJGiEa
zRFehUdIsxNeP7xcjDigSeSVbWbHHvAuCJAI0LKO24mOUh75JKwSTLiSe/5t+4FAwZpv5XtbOGRM
HskUJuZyPwZMoM4+X+4y2qNzoNB7V1HAvzxRix7pTLxz1V3odYnA+9LEOvzV5c4GaeOGNUZH+9rj
+9kaOqU0d+jOAINzbouoUoKSmUSfsRBHYufHRg17WFMDxxkfOfWnoxFhO7CN9/NX+rNvMVVWAxkm
51/0SPcGJI7ryx7LNG221dt5suxKEEDkIu7U/wXjCkj9cpKKnrE2anZjkA0vWv26IbBkStJzjBzc
AWHGt0HlKGqYhJJ00dw/hdgpqSSMlvVOBwMrb7FVsP/2wM/12dnJSFiKAOHckuChrpU8cE4q3z68
Lygzn+TketZEd0OZqsWoCqtcXhVi5MOcxygEl9BejbPd5fOH5CPTJewwzpAkq6jBwS1YXC2+rXck
vegCuS91rsNSMe6/db+1PUN6ibggm6irnhWsjarmFirpdDkqvdyTQ3rFQXKZvNIgVOH8XqyHWwWc
slN3D6nc03P9CTkYt0mFMADz171FUhGUhwcdWXjK0pj4yh+tL4q+dLrtE199+Y68KVI6w0pDaPCJ
50E4ygTzISkpbL6lEZuGLKtlgyv7a/WWKJkK6OKsYasdLV/bz34j/jggJcD69jJ/pYYj31YnSTOC
NMwVg4hJe07zRU+5GWv3ir/fjtdNaBgAXAO23bacgD/iq3mxXBInXv2zWDf9QdWtEUfxEWWUcEh5
ftSjTIhuwgUphBSCKod1G53LsJOFe9KLafd/z/D/PhlFsv22RHeObERmPTFttFGFjnCMfZ6g5s/Y
OIVJLHoaoRbd/03SmQXVk/Brbr5s13rmEh8uhKKfXsix7nDLufGddO1oYX4+9evURAC7gAisXPFL
1+PWtU8oIfW1oDa2w4o3F2Ki1FFZRa9mh+f1E+PIDy41UEZtL6l6PLE8fQkxmblJ5vCshQwLtmj1
WSRDdKI5fFD9UwXFu7lF9Rwp5IAqVVabGBUvWcLca49vNYTeH0OEdOY9dkRJs8keAXtGzp0M3C9/
Vh4PyWL+A55TtR6c/LmKpU6isBvzwSCJNzr+miERBvPMk2ali7NaAb5ha6i1ehcZW7gXBpBrR7JR
OrtjVz/U6TptteA80UhoMvbg4yfdyot7j/b4rS32PHFluZT2SxqS2ve1o+PkM1nwsZdnXOd2hViX
xJ12U2VfwY6ELEDLrjUHTubA6yaSqkNngPbYF2q7uIYyVDSNtmGjYmGpUgGCdvzK9IiM5DnFjIgU
jwF+1cVuVV8SQk7lttieYeAkcGIkXIBWY5k8QY5E2Kdr5rPVn3k/8n00ZCz7Xvl9GWca15HB4MRo
euKPma7s2e1u6QNul8MaVzdvn7MZRnk+PvG2okTVb9cj6UVaEIGm+QOkNiLzrQiGNKMHXg/Ovi/h
raclb5rSxZB3eTykWlQMU3U7b9JOIRLbTaKrtmhW7oOQmkkbBQM6nlMtT8j08L4hSOC4oh1oo2BE
rtYtfub+y/O7cfqKUK1ODRNCNupbPJcCFdBwbOp5u3PLi/p+xHlFwAMSeM95MC0MlQyk5t1Uj/ep
g0lyjpHGdgBTJMkGf6DyJzDIYKUGiKl5vcxeNG4Y8/Jpj3PTxmnDA0qrVw3oJhUnpuiJwSWMUoVX
ITmAS0lIXIRp05HsGEToxKmq5px5e2q6CsyFK0LrL3ftoY72z1+kxgmNCHtp6Ykst1FxtqXCf+qG
KFnbGjFBlZVeeDqknCD+Qk+bYlC/tJVwXF9ff+L/maQ6zkuc9Ng1+PAimqz7nnQS+/f1Sj/A5wPk
rAJvDf2JhOaOqTY+XYeTfgPqVLHF7vdnvR40BcEJjVnQkF6b5tzpAQ3SjmDqdtBrgjzYsrlIuJZq
90RCiY2C5Us7Agn+/A5T6DBkE9Jiiqh2taZ+loPSHJlEJaNZZkXKZarDwY6s4flPXctkTKcqZ/x9
0oEgiviqU7j1k/00FxV0O//Iw/qUTwsnQBDlYqgTWADnoQ34KooHVbeIw43+g4LunTuLCzlmdfoz
/tpBRmLHbuy+7/OFS3Yj+tQWC87iOnk3Kq9qQjGBf9a9grt8Baw4UAkPNQxv42Eb/3270kZPQKFj
87gwb4jnaTt85E/fwuuIEjg6dl/TR3NYsraKbBo4/nMR9MUAcPPqngWTIk4Wt4QFPPnBj7V3ri2c
JzUx/AmriKcNuWNvXS+ZiDjqsa2xOeA6KoVKGVlT3FKJVccXPb0ic8DDmIu2kSJNMvBEpdJTmb57
GAaxHMDGEPR3M5icYdz9p07H+dhGMNb4AqzmFFr5ZRBPxtmI4i7HsnP9e6vs4avRJ0X8YS8/CZ2d
mp9Ve+tpLPOUhadR3B2LkPc/D1ymZLEezer5AuCEcZ/35sAb5GkSkrWgIHBqDnsI+XG9TcL+Ptr+
rN49YlXIrbkvMEKX7CzfU/RRxyFjLsYBeVXaE4IeQx3oZQMluOx641Y83Qd7+FaJwvn9QPYbEb1b
qaE9X44M8r3a3HIRttfqthA17dhO+/b3v02LCmVLEAPERVGZn3ETpEO87vDziK1FCfqDpddkdoeD
r05IkfhDqkpKIBpfkllRddUX7aJ1/omMEiBND5gGXzydHBa5OS2HMYctCFbi0LQDZ4gsATZ9PEdC
NZN786x7QE5ERu6YZnxqT6/IL1UDn3rtxA8F4t3v/UwG/Iy9PC9bQ+qMaC7SvTEC+Wlbg6UW0XFr
fvjFXfbEdNbykvm4tQEKnLMb8TzQrIaOPFTGldsm12HDhz1R80prsXYl6CMqGK8uxND/4MK2oHft
YunnHcwd8+FrPSb7XvOdiu0sIGjldwWW9qPegclvQkYy82lP4CgZiilOzaBTqCo3LSJPMYh6dXu5
u+IQ8eSrMilCW9qQrBcYjyfGP7CesgzbKFC01+CQr2DxXQMj/awH+SCy+AIh9GRMJNDmJBQmZ/6b
86snYYhSgH3C4Bcc3O8Qy1f+I3sa+E6r+w9HIFeoU77Mb6MiD54dSR6fZ7aFsTvubtGirgW2PX1q
sGiEGuO6QzeOmcrpXrQjjxx9vVFd6Vw/zIXGcxefF7PSPED0npjK0NMw4YW+4hfese+b8qjYrPKG
HerfFAsD0qqWLI+VTVCT9T7aaCPFKyZ1XE2HB6NB58J0Xa5O2nun3GnIV1KBKh3cdCb7JFxOzFau
HOlwMjYULetwWa6cCm3rDDsp2g9EmvBOFEs++TQSRh7qO7tjtKPr9wQTJpzzc2Ht2pZWQ/9qfFSD
HF9PnZM/uO0JvbnhKIn86E0bgXqle63+WCUlbigbOOc2Xf4/ADYxdHr6kzCMQJlUHPXgcTGneVeV
LeUwfPAxNiibm/lbZ/jDEXUK0BvjYzDfbgf71BDKUMJjKfzRDtJdyZp6TJZr+D739oORnagGL6CV
8Ieot1ACLaHBeBGv7tiJJe8P5kskYzM1CPF4XvTVc8vcS6Qb9F0ONhG0x3K/bJnpe/DyAt1z9Duk
bvf4t+vroOzPYKoeb5p7+EQlHN6CSj1WdzXCqEU+5q3KgRL5TZIg+Cif9atvNgT6ygldk4K7ED/w
zN8eDWs0SEYQDbBKucIys7+YDgMgZEDwtmubtBQBNwBYLTi5Z+MXzQKXMHQaUTfm8lFOMojGsh1S
fhYSADzJWYTWfMmL8IIf9J0nl5QKjGHcI8Vu3tDZEW6vJLSCJ0rRuqUQ4nvqLy1URuJJd0n797I3
Csha8iy3rt9VLLiTibJmUXv70I0U3yiEgUZx2mRL4hm5FOzzhdo6urr756pL2qzB/eYZ4mfjpe8Y
MvZP1QsJ2u7uLrFn8MohS8Sq4EBBh6mBjpNP5SdkNLxsFvNgOAwBkBxzNu9h7HBMTpTcwy34eurP
/QWIoioiSD+Z4PJpvjMi1e4eYmBcHrwJvM2GtTMzfjdbBnXGcv8K58H0I8VIavUqwen8qGq0CkIW
8jBBzM4M6js6kBfgGUIobLvMsS8eNQh1loDvlQK/N2oE6WJfWmdOg3TEa2IBXa517cFV1mnehyO0
DhBUJMFpkG0VGAB2IAsquEPaBM6jdpCGsp4q990zqlca1WagqBhkyjtyIpDwuKXBQjzdk9rHGqoX
83dz623talOiYH1M+gReTiKNGlfEKwZkBSFWmtcmbhmS+dI+AZbAQDBg9KlIYD5e59hcbnlBJOJt
c6f8cnmbC+jQrl8GvjKW4XsK/q8mauU8rzII4cp+Xq53McaoZwsxw0EUFY+hr7s2ZWDdKJ/c23SN
ECU2eyOayJ+dBPk0bhaPKzSnk1sQHvAQ19s3vNknvdO2y1ggjc1pQ9v3EJsVeBWLsTPD3b5bDoSo
kucbbUj+aWuUwBIwJalVZrGCJFzdyID1N6M6d89gBeusbfGGJicIDXmaHn5W0pKyGSA3UrbXLyxd
TXEYw53yFatFKGN6Ckl3fQDWU9g5vDBu6ScTy+AMM2EdMVHrdTQZBDit3JxcirBEjXMS7Ug75+8c
KgC1GVLdTj5sZ072WC/1RfGo6aKS514DRRf0cfWCI39A74lQCFWYevI/p6FjgntZnST8lVghSl6x
kB3I4c52FZ35GkyaDhZALCu6Tm6vqBfPpoYiYwi06wzDfD/6Mb7OppZVNAOYXkMjrps1PwvnBAN4
NzSQwEwveiG9y6ouAnggLtu9OymgpeuDDAEDu3KaTsjsElixyMX6v1Oj+zZDpVubq7e7TrY0tmtd
1ZYFiHPYkV3JCnA7AyLbCHa+90KR/I8utsNmvokPguWN1Nv1zRVV6wn4VydG5/BiI6S+P/pyeIe/
jrn8OxW4Er2kMptmSBvfw0YVD3Hi3/+JDEV0KR+LRPrt5VorsMyheb5yaAlDcge9XaeMjxO4UpoZ
4Uc157VPgJoPwrlXR1IHONLhWLu374rNSVkWImkQkiFKRvk7x+Y3gpWTsOq/U1ECxNSbzj+frX3q
L7bJpNKSvwa6TtM+FfiTEErE8WvJ9JGLpLeV4ex37V7J0XjPjrTY0dw8ZGMzIrjy5vbPbSqDFgTE
LR+z5/vMlmwDgAAD/tzO9nzUbL7Gp0K4uAHiOcXJ6IFei0XfbXzCaTmiibJ5Os/jZFMXI0IrEQ03
XRWWexspnqg9DXQCBcpNhT98AmIH1noHaaP+vFYmtUzoKtJ2jap4G0oNUAhvUFlWqxeJSDSK29/V
YaqXqXJRLAv7ct33PJL8we0Dc+wzrw+qsG1eoeHdOZ/d3bldlJPr3O60e55r+eJ+SlR1wRy0IpZR
QlMf/erTRb/22ELdF/mOeE4vvMiCzh5a1lOzywLB36VBgEV8wZlaZOsUn99j9Tnp+VP/rVOhwI7q
u+AgMd5pde2Wzkc8HFw0xKLRJh1vuzK5pGZ4GjVyiaCCwZYnOC4wrYMCuafDExN5FlVEQ/1ZpbKl
WDfpnKZqLBf/wgJEX2etSoEkynm0cfC0RE2xafX4uyBvijgRqJcUModpJ2A2TAoZ/jppzBGmOh+i
P4EB+YkLo4ymdmq33aBEYvYfSnP3bFrq/0UcrMfatTx+wXgJzzJB1R0xVX48HuCSbrqv25u5krqw
kDltpfqQS5HxuZ5VROyfyHwWUHiFRPOhAMMvP87Hs4aU8WStGVZnIcZA+z8xkVXrGS+Dc+tomJ7a
zXINYrzWbmiExkD9JLQmvu2a/noPre+pTIhb3F74uOrNhfCmMzfDXTUtUKh6NGDe8SX8p7s8OIiW
BOx3927vkA5B11XNhlWN3sXhiFWqMrBg9rgN0kl6gsGwXi4tUPI45P/ZBDAEhenW7dZUrX6KRgyN
cm/698z2PcbEp+733d30GrBoY5c6qTvVXL3d0TeVNXIWJEGFMwjgXYCtk9ItHlsPxecN/BFBFJ2A
kvAzEMBdFDNWStVUmlzqNZUi53G8qLUgh3nwX2iAVLoB0LdX7RGe1i2h7QKByqDf4f58fQ+yuA9S
w3z6IpQGvcej7PExuFPUi7+xZbFeWURa5J8ox1p6u9RNkCXpESiAAD3yMRsFJuRmpF0kNBpZJuWd
OQg0gs+7N1sf8t9gakWRzIQ+IrnR8Eu7dlC8KK1YKFc1gbP4rWDbPOD512/fFmRiAhcD4Od4UppM
RSf2EplL6qDseZtGisbX03JbiqaqQJH+Qr469USCcy0/uATLgl4dxi7zedjmiJtr6E6A0bDi4RKq
zDhfLuhqDw2cL8TD8Pw3ByQtxtu8wVBH4WZbMI685et9vO9HqDR+yLKRJyTQogJGU8oZPpSJQg8C
1ah6oU6w4jbfbkOaeHvTeWLe+634+6MtVpQOCGKcLqN75Oy1w6JIlqS/7mcmd1z9w9X3d1WXZCX8
PjT90VZHBzHaf9URVZraRpLE3ZD4f/7WigkWWi1u7ybONiPLbJJHyzuFVnI3p3EgArjSulD+9dBR
PjRIeUhQ/B2VM7iQraw3/WCbowTBeEQZsOgFXutEKkRgF25H6RazAL2oqQoLA+3sDI3/03ZbhrDN
CdreMdl+KoqkmN4kTgpBthqMwX8soa24WVwAS3rrEgVe1A+IlFt88t6vb8Lbp2P2qlEGK0avqpC0
FiwYT+FFbeYUHfSpQ2ZmST3K+VvmpLoVruGKOY99pLQ+hr8pKim4Zbun70FryxnlQySx5M+I1i6V
sN4jy5j44DCK4c41UPtavs4Bn3zuBnnL8E8aS1HC3qE/yl0hauhHtNFS82RFC693IroNR5s10Chr
HVccJo41SyEgYXqQ4/bxxRT6wLumiAnW4G4SKKz7a4YUyuj1oO+psRA6PYBzMO7qubrojm6DWzJ+
3LU9dMNw12RgGY+i2OjnBBHAfywxKN0hJrin4saeJ0P7tWaortHQaZiBWkoO2hShqnI2yl1kkbKk
G1W8rz8lvhq+OyKKa+izkuCeKkRMm4rqLlHEXxNSuCO7o6ut8j8g0kBdc8xhuVLvf39w955nRABl
jau/JuwtKuVWJQNFJfJhJX+R1bm6fzA+V5OTs/chmUP1GoJKUfsf/dBMUoWc3dcVn9eIuOkNUE0I
Au97fOSv864O1bsRCrKKBTEg1aMA37xg6BKR7O68K+IriDODPvp/y/9+3HcTtA4UsPdMGJpf1oOU
YNfFzpD+K82iInh80XQZSuTodA8t6elDKcjwBO8bp3JMGvZdbQjCoA/tsoCTTD1slWUZTuAQCh6S
Hu1P43ymhaulefCmtJXaFbjhtwSbDtDPxlG6v+1Cnz7WLSukCUTCpM4+b8WzjYsB7SioySwMIG59
qLWyIzMjmxURXoDzC4XWePGBaf8TwWM6jH7a9ACrUSWv7/Ob0ors3m4rZh41LthJy5K9EAIigXIY
3CysotLIt3PxQ9XUUbx7e1nR/AorRazSk4X8forKIu62Rk6e3dtCkEa6byqbBC5red2RC/C3YVHk
JafVz6Dtrkj+rg/V0nmdPDC9NZFY1r7n1Cr7Awbd6lmSBXnMZW3Tqf14y53lfZKKsCtdUb1okkbM
SuMG47jJ/YhY3KpmblL7uxppz5jojeBccdNAopGwQuoB0Y2GIhSt1NAX0lTBz/Oo+cqGFFTvDsKl
4/35eUcUwhn2XXo/NCzQR4OWs7VyS0/abS5FMc3aE01qs8znvExGW6NeLWBzYUPT0LyhWHOoVlBa
Qf2ZC1v68luYfpaMWJiLJN9SFnedaIuHO6hKTNyKfWqNNOySc25bAe6dE9GrjLHLPoI41ow3Tl4x
b6SS6SaYcsuH3i4SltJU28aggOc57dkhLm12Q34wHGKK8Slmtpt4CFzY+GPO2atvKA2UE0LJRH7L
M6ZAmeuWm3ejPglk4AsWiOZekRfht1Zg00EN4sD+X0zU89Jpw39AAUmzkJu4GUHo/h8RvWgWUJ45
4rj8t6W4lzsFZ/q6yE7OIA+i+6Hcm7j/OLTzFJrdQ8abpTaUl2gnogANRwUc95D4l+Slie8hPtt0
x07/CUPm1bOdxhEt52SCeFVmp/B1IvfOqJiKj9dND2jeDlAX1jaVTOTcSYVIRmdQFaw4XEhIeX1h
hZQR246N8wiP6zHwYU6h+zI+G0OmCfCKK3cFXHCd7D+QyAZUjgTNCl5tWf4Hg6sHXyHlQzfBGFBf
NmT8O8noBj5FXPbPQ65vPdRVUoipLgMRrlLTFFWfMy8YAQQc4xxXk0UHkKhWgPdaouShV/ZcDAwt
E9Yfwkinx1Cz2GrSLJyGvP3DDxokpwhFG3NTHBTSmx0gMlDHW/jqmAleokE34/kCY5Ylqbg2OkPg
x/9etyDbq3yOF6RFwSY3UA/Hx9DXg/sH1S7ZYHz5BIypptvcERnWzn2np7eMMgv/k75fXHVen/UZ
l6FDRa1Gb/IgjLcIr+BFAn5qIFZZIpOfSsmthqoxCj6o/dVNAMkVZv0w8XvH6H0Oe6qo6CRlqzUD
V0V4jEF0jeUPg0zNAEEtZ5UH5VARLAF8BQm2jtBhZVawrdveH96d+aER1fdLQe4cN2FDASVfOyeB
m4XlwgIahg5NM+OTZsfFMQk7RN2ThzZFEXfaA+D+iOb9D1d2HQwmy4fObViddBEYVF0HjuSlucDo
tDjMqejlfDuwLtlLA8kqXM0tnY7RFi1B8tY9yFg1DK/qdafEJnCCbeIsT0Yh9Ufw4Tmyei7USsZF
pU8xTaIa7qN+fKtniQBJhxzyHR8QESVspvnl1y46Q4mqhJg379OqaQJUFsOtB3Y+qV6nBwcwus46
j87gJ9dOtT2o72mGHu6k5Bm8tgQ3h7I/9G5HZ/RYig2UMgg6kyW7debAwknH9OABjHVsCuU4Rdqd
OiPCGxNDk58BXW2FYgKqvPRTYlaa8TEsUm4hKGT1Rm0oAXwjePM4m9zYgsL6prtyneLr0IgFmrhr
aT+CZjVccgpqI8U25/N8YPbhH5bXlMSBtAjI1ILd6siwMX0bUhcpEb5pEbrVyCTn/ZWbtyQIdsBq
4BycANgKZfkauS2nJPAOYdsG6+/j61w69T2HwfhtdFRoLZFFwQqzs0jnpUQRbOKV3mXml+wg98LC
Z7ES5FhKHHYl90iRTZkZc/qScGvqZCytBQOp7Jee7pdd4ZI9psu8wUGP2jKAllVuC7lqufwCvnTq
R8xdfgEweYRWiXPETOsC5yvjyC7mggE2KbNCIsRB1mDg6p/LOiaJ/4lxDIkiLdRzErlN0T2Exbxb
fCLFLikneVCBUTsfpzu73Y5yIl2mR8YUh7L5RXD4XnkvKKD1PNdBifItzFnF0bGRdWi8x6ww30Xo
CHuSwh54wMaGsf9oUfZEhCc4ecapUwuwj3LUfALwwbnF1dEe5BNCvSNakAx2MUEQdhE1e6nJMz69
bOt8QUxGgJCkED42kX34KwR7SYFdLZzRHnTt1g7DDETvKVRpMyaiDPuI7AHCGQyqir2uxKuy5omF
30em9+IuEoyXyAEywljpC4lEe0BZ6K7MY4cHu1rAXWWOrqeHPmmGSt+n5jT2ueLFuTh6PdBXp1Nj
KD5mia0jIH8WSZpUj/glCCtt+3iyMV9h6iGILtfgssy3lWOEUQZnqKxvb6YvuVNPJwLYpto9AitV
EZz2Ar0J8WxLCMwQmwGUudqEwvrxr8eg5LohUiO3iKYlI6YKJ5O4pSzk2f0dRc/13dZR45mj+L9U
32fWIiiGlwJ4VlNF2v2TAwFTc2zsmnOQBpFP+Fe1QfLNd/8VLmxjAC++54T9Pr6LMj30FahJ+Q0m
IWsadP2F1+eiIlwWjPU8baA3Y7TbcbomBDrISoEwVfJWaqQMbZvHggBKczYbPRlpdwXb698iZ304
QFHMHk7U1zIwO4FpXDKD2RpPQiPMWvwpks+bQhILgvrcB4RLyHDozWmiBRpKzjasWV4r+CB8+3AC
YXSNC3a69jiLOW1rT1MfjCu1J+Uk9knFahEMtig7F4CmWJVdnbNo2VaDQelWKtKhVJo2Ubh/q5VY
ULO9aYrfNtbcNFaxYSzLVyUrNEsELYU08y03rAHVuDAJnZx2i7Gyj8qc9wqjfUQ+Sqvb7CZCerp1
+EVS9TbsN4IKkoBGM2Tp/fVrpbqVEFUmBa6gFt8d83lbi7LZ3ZboGTd3HgeTsS94hXgDAwfmYkJF
uxtmUos4Td6BM028xcfw3n12vhUADJPeUvQk70ZnNtMQ3eIEyV6zg9b244ILQN4Tn+NO/aWvfO+I
CZBsby7HD4/GRBceitDOcoq0EKegFqvbo3xatbs7cMN6ZdysKtbDni/hxThtwlqTR5SNMpaUKXot
Hyqm8kO3BzWt/R9xX3GEL82ds6ID5tKWo04rSYICyPvArY2tLE94UncAP5xTXvNO4ap1hrplUjRi
BPhCZN4MgdTnMv5Rrhc8mbQKuqOtyL0tt0ktGNpaugrC/Z1Ci4aKTJ+R/B2KNTxiqt30XAlReAKS
1Ka5NT5Eh7doQm9OkQ10ASM2gwzFUUBMawgSWzHQmWbzV0DRqNGyetV1FtI33YQrBmb0rrQ2gBk7
oXfMfMMkpJVKa775jeqpk6ANR9QQj/Zf/vApyk5Q9UczNbChqiWLL6fiCm9hI/MlLC+CwRF46rUD
bNKYrB8LMYepRnwQ4qE4+oMpDa1PGivyqBjG/bnm3NDeLsvWNMlOoQ6tgfudp5mEAMNAozw3GLX0
o8Krvn6YBgkXCgJ2cAlXlJz8p6J5KqKZeRbBMyDo4KoUT3nVOOMmWI3xC3dAQKsWgqu78tifbkpn
VE2CWtdQwutu24y7uTI9WZaelSxwg3aoRwZyiy0ya/pR8yMCORp/phkb4Gb1Yve8R2U+dxNAtqYy
a4E4Rk3gDkqgwGVFNg3EI5QiYd2trusP+cf14qaiVZmDQ86u83MPAZek2zwc2UF1DAHBzCO8F5Ku
7M92RYKn8clTfDC+sUYjOq7T7AxKmHTcBzII9en2GI318PLxjnELJD4pJYf+EUKbM5YV5iBTyGLZ
vG/9LzPTsFxFazm0scyzRPUvNit7fsi6IqymfZ4ajwpBmxpQoRsnJSKxMZg96mT8397uTIsb/AU=
`pragma protect end_protected
